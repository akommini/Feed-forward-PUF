** Generated for: hspiceD
** Generated on: Nov 25 20:52:11 2014
** Design library name: Project_658
** Design cell name: 64stage_FF_PUF
** Design view name: schematic


.TEMP 25.0
.OPTION
+    ARTIST=2
+    INGOLD=2
+    PARHIER=LOCAL
+    PSF=2

** Library name: Project_658
** Cell name: Arbiter
** View name: schematic
.subckt Arbiter d1 d2 q vdd vss
m12 _net0 _net1 vss vss nmos L=40e-9 W=90e-9
m5 q out vss vss nmos L=40e-9 W=90e-9
m3 net5 d2 vss vss nmos L=40e-9 W=90e-9
m2 _net1 out net5 vss nmos L=40e-9 W=90e-9
m1 net4 d1 vss vss nmos L=40e-9 W=90e-9
m0 out _net1 net4 vss nmos L=40e-9 W=90e-9
m11 _net0 _net1 vdd vdd nmos L=40e-9 W=180e-9
m10 q out vdd vdd nmos L=40e-9 W=180e-9
m9 _net1 out vdd vdd nmos L=40e-9 W=180e-9
m8 _net1 d2 vdd vdd nmos L=40e-9 W=180e-9
m7 out _net1 vdd vdd nmos L=40e-9 W=180e-9
m6 out d1 vdd vdd nmos L=40e-9 W=180e-9
.ends Arbiter
** End of subcircuit definition.

** Library name: Project_658
** Cell name: 64stage_FF_PUF
** View name: schematic
m2096 net04309 net04302 vdd vdd nmos L=40e-9 W=180e-9
m2095 net04309 net03543 vdd vdd nmos L=40e-9 W=180e-9
m2094 net04489 net04483 vdd vdd nmos L=40e-9 W=180e-9
m2093 net04489 net04482 vdd vdd nmos L=40e-9 W=180e-9
m2092 net04519 net04512 vdd vdd nmos L=40e-9 W=180e-9
m2091 net04519 net04513 vdd vdd nmos L=40e-9 W=180e-9
m2090 net04459 net04453 vdd vdd nmos L=40e-9 W=180e-9
m2089 net04459 net04452 vdd vdd nmos L=40e-9 W=180e-9
m2088 net04429 net04423 vdd vdd nmos L=40e-9 W=180e-9
m2087 net04429 net04422 vdd vdd nmos L=40e-9 W=180e-9
m2086 net04399 net04393 vdd vdd nmos L=40e-9 W=180e-9
m2085 net04399 net04392 vdd vdd nmos L=40e-9 W=180e-9
m2084 net04369 net04363 vdd vdd nmos L=40e-9 W=180e-9
m2083 net04369 net04362 vdd vdd nmos L=40e-9 W=180e-9
m2082 net04339 net04333 vdd vdd nmos L=40e-9 W=180e-9
m2081 net04339 net04332 vdd vdd nmos L=40e-9 W=180e-9
m2080 net04302 c57 vdd vdd nmos L=40e-9 W=180e-9
m2079 net04482 c63 vdd vdd nmos L=40e-9 W=180e-9
m2078 net04512 c64 vdd vdd nmos L=40e-9 W=180e-9
m2077 net04452 c62 vdd vdd nmos L=40e-9 W=180e-9
m2076 net04422 c61 vdd vdd nmos L=40e-9 W=180e-9
m2075 net04392 c60 vdd vdd nmos L=40e-9 W=180e-9
m2074 net04362 c59 vdd vdd nmos L=40e-9 W=180e-9
m2073 net04332 c58 vdd vdd nmos L=40e-9 W=180e-9
m2055 net04333 net04309 vdd vdd nmos L=40e-9 W=180e-9
m2054 net04333 net04311 vdd vdd nmos L=40e-9 W=180e-9
m2051 net04513 net04491 vdd vdd nmos L=40e-9 W=180e-9
m2050 net04513 net04489 vdd vdd nmos L=40e-9 W=180e-9
m2046 net04550 net04521 vdd vdd nmos L=40e-9 W=180e-9
m2045 net04550 net04519 vdd vdd nmos L=40e-9 W=180e-9
m2042 net04483 net04461 vdd vdd nmos L=40e-9 W=180e-9
m2041 net04483 net04459 vdd vdd nmos L=40e-9 W=180e-9
m2040 net04453 net04431 vdd vdd nmos L=40e-9 W=180e-9
m2039 net04453 net04429 vdd vdd nmos L=40e-9 W=180e-9
m2038 net04423 net04401 vdd vdd nmos L=40e-9 W=180e-9
m2037 net04423 net04399 vdd vdd nmos L=40e-9 W=180e-9
m2036 net04393 net04371 vdd vdd nmos L=40e-9 W=180e-9
m2035 net04393 net04369 vdd vdd nmos L=40e-9 W=180e-9
m2034 net04363 net04341 vdd vdd nmos L=40e-9 W=180e-9
m2033 net04363 net04339 vdd vdd nmos L=40e-9 W=180e-9
m2021 net04311 net08593 vdd vdd nmos L=40e-9 W=180e-9
m2020 net04311 c57 vdd vdd nmos L=40e-9 W=180e-9
m2014 net04491 net04467 vdd vdd nmos L=40e-9 W=180e-9
m2013 net04491 c63 vdd vdd nmos L=40e-9 W=180e-9
m2012 net04521 net04497 vdd vdd nmos L=40e-9 W=180e-9
m2011 net04521 c64 vdd vdd nmos L=40e-9 W=180e-9
m2010 net04461 net04437 vdd vdd nmos L=40e-9 W=180e-9
m2009 net04461 c62 vdd vdd nmos L=40e-9 W=180e-9
m2008 net04431 net04407 vdd vdd nmos L=40e-9 W=180e-9
m2007 net04431 c61 vdd vdd nmos L=40e-9 W=180e-9
m2006 net04401 net04377 vdd vdd nmos L=40e-9 W=180e-9
m2005 net04401 c60 vdd vdd nmos L=40e-9 W=180e-9
m2004 net04371 net04347 vdd vdd nmos L=40e-9 W=180e-9
m2003 net04371 c59 vdd vdd nmos L=40e-9 W=180e-9
m2002 net04341 net04317 vdd vdd nmos L=40e-9 W=180e-9
m2001 net04341 c58 vdd vdd nmos L=40e-9 W=180e-9
m1984 net04305 net08593 vdd vdd nmos L=40e-9 W=180e-9
m1983 net04305 net04299 vdd vdd nmos L=40e-9 W=180e-9
m1982 net04485 net04479 vdd vdd nmos L=40e-9 W=180e-9
m1981 net04485 net04467 vdd vdd nmos L=40e-9 W=180e-9
m1980 net04515 net04497 vdd vdd nmos L=40e-9 W=180e-9
m1979 net04515 net04509 vdd vdd nmos L=40e-9 W=180e-9
m1978 net04395 net04389 vdd vdd nmos L=40e-9 W=180e-9
m1977 net04395 net04377 vdd vdd nmos L=40e-9 W=180e-9
m1976 net04425 net04407 vdd vdd nmos L=40e-9 W=180e-9
m1975 net04425 net04419 vdd vdd nmos L=40e-9 W=180e-9
m1974 net04455 net04449 vdd vdd nmos L=40e-9 W=180e-9
m1973 net04455 net04437 vdd vdd nmos L=40e-9 W=180e-9
m1972 net04335 net04317 vdd vdd nmos L=40e-9 W=180e-9
m1971 net04335 net04329 vdd vdd nmos L=40e-9 W=180e-9
m1970 net04365 net04347 vdd vdd nmos L=40e-9 W=180e-9
m1969 net04365 net04359 vdd vdd nmos L=40e-9 W=180e-9
m1968 net04299 c57 vdd vdd nmos L=40e-9 W=180e-9
m1967 net04479 c63 vdd vdd nmos L=40e-9 W=180e-9
m1966 net04509 c64 vdd vdd nmos L=40e-9 W=180e-9
m1965 net04389 c60 vdd vdd nmos L=40e-9 W=180e-9
m1964 net04419 c61 vdd vdd nmos L=40e-9 W=180e-9
m1963 net04449 c62 vdd vdd nmos L=40e-9 W=180e-9
m1962 net04329 c58 vdd vdd nmos L=40e-9 W=180e-9
m1961 net04359 c59 vdd vdd nmos L=40e-9 W=180e-9
m1943 net04317 net04307 vdd vdd nmos L=40e-9 W=180e-9
m1942 net04317 net04305 vdd vdd nmos L=40e-9 W=180e-9
m1936 net04497 net04485 vdd vdd nmos L=40e-9 W=180e-9
m1935 net04497 net04487 vdd vdd nmos L=40e-9 W=180e-9
m1934 net04530 net04515 vdd vdd nmos L=40e-9 W=180e-9
m1933 net04530 net04517 vdd vdd nmos L=40e-9 W=180e-9
m1930 net04407 net04395 vdd vdd nmos L=40e-9 W=180e-9
m1929 net04407 net04397 vdd vdd nmos L=40e-9 W=180e-9
m1928 net04437 net04427 vdd vdd nmos L=40e-9 W=180e-9
m1927 net04437 net04425 vdd vdd nmos L=40e-9 W=180e-9
m1926 net04467 net04455 vdd vdd nmos L=40e-9 W=180e-9
m1925 net04467 net04457 vdd vdd nmos L=40e-9 W=180e-9
m1924 net04347 net04337 vdd vdd nmos L=40e-9 W=180e-9
m1923 net04347 net04335 vdd vdd nmos L=40e-9 W=180e-9
m1922 net04377 net04367 vdd vdd nmos L=40e-9 W=180e-9
m1921 net04377 net04365 vdd vdd nmos L=40e-9 W=180e-9
m1909 net04307 net03543 vdd vdd nmos L=40e-9 W=180e-9
m1908 net04307 c57 vdd vdd nmos L=40e-9 W=180e-9
m1902 net04487 c63 vdd vdd nmos L=40e-9 W=180e-9
m1901 net04487 net04483 vdd vdd nmos L=40e-9 W=180e-9
m1900 net04517 net04513 vdd vdd nmos L=40e-9 W=180e-9
m1899 net04517 c64 vdd vdd nmos L=40e-9 W=180e-9
m1898 net04397 c60 vdd vdd nmos L=40e-9 W=180e-9
m1897 net04397 net04393 vdd vdd nmos L=40e-9 W=180e-9
m1896 net04427 net04423 vdd vdd nmos L=40e-9 W=180e-9
m1895 net04427 c61 vdd vdd nmos L=40e-9 W=180e-9
m1894 net04457 c62 vdd vdd nmos L=40e-9 W=180e-9
m1893 net04457 net04453 vdd vdd nmos L=40e-9 W=180e-9
m1892 net04337 net04333 vdd vdd nmos L=40e-9 W=180e-9
m1891 net04337 c58 vdd vdd nmos L=40e-9 W=180e-9
m1890 net04367 net04363 vdd vdd nmos L=40e-9 W=180e-9
m1889 net04367 c59 vdd vdd nmos L=40e-9 W=180e-9
m1872 net03549 net04550 vdd vdd nmos L=40e-9 W=180e-9
m1871 net03549 net03542 vdd vdd nmos L=40e-9 W=180e-9
m1870 net03542 net05098 vdd vdd nmos L=40e-9 W=180e-9
m1866 net03559 net03551 vdd vdd nmos L=40e-9 W=180e-9
m1865 net03559 net03549 vdd vdd nmos L=40e-9 W=180e-9
m1862 net03551 net04530 vdd vdd nmos L=40e-9 W=180e-9
m1861 net03551 net05098 vdd vdd nmos L=40e-9 W=180e-9
m1858 net03545 net04530 vdd vdd nmos L=40e-9 W=180e-9
m1857 net03545 net03539 vdd vdd nmos L=40e-9 W=180e-9
m1856 net03539 net05098 vdd vdd nmos L=40e-9 W=180e-9
m1852 net03557 net03547 vdd vdd nmos L=40e-9 W=180e-9
m1851 net03557 net03545 vdd vdd nmos L=40e-9 W=180e-9
m1848 net03547 net04550 vdd vdd nmos L=40e-9 W=180e-9
m1847 net03547 net05098 vdd vdd nmos L=40e-9 W=180e-9
m1844 net08551 net08545 vdd vdd nmos L=40e-9 W=180e-9
m1843 net08582 net08575 vdd vdd nmos L=40e-9 W=180e-9
m1842 net08582 net08576 vdd vdd nmos L=40e-9 W=180e-9
m1841 net08551 net08544 vdd vdd nmos L=40e-9 W=180e-9
m1840 net08575 net08884 vdd vdd nmos L=40e-9 W=180e-9
m1839 net08544 c56 vdd vdd nmos L=40e-9 W=180e-9
m1832 net08576 net08551 vdd vdd nmos L=40e-9 W=180e-9
m1831 net08576 net08553 vdd vdd nmos L=40e-9 W=180e-9
m1830 net03543 net08582 vdd vdd nmos L=40e-9 W=180e-9
m1829 net03543 net08584 vdd vdd nmos L=40e-9 W=180e-9
m1826 net08270 net08264 vdd vdd nmos L=40e-9 W=180e-9
m1825 net08332 net08326 vdd vdd nmos L=40e-9 W=180e-9
m1824 net08301 net08295 vdd vdd nmos L=40e-9 W=180e-9
m1823 net08301 net08294 vdd vdd nmos L=40e-9 W=180e-9
m1822 net08332 net08325 vdd vdd nmos L=40e-9 W=180e-9
m1821 net08270 net08263 vdd vdd nmos L=40e-9 W=180e-9
m1820 net08115 net08109 vdd vdd nmos L=40e-9 W=180e-9
m1819 net08115 net08108 vdd vdd nmos L=40e-9 W=180e-9
m1818 net08146 net08140 vdd vdd nmos L=40e-9 W=180e-9
m1817 net08146 net08139 vdd vdd nmos L=40e-9 W=180e-9
m1816 net08177 net08170 vdd vdd nmos L=40e-9 W=180e-9
m1815 net08177 net08171 vdd vdd nmos L=40e-9 W=180e-9
m1814 net08239 net08233 vdd vdd nmos L=40e-9 W=180e-9
m1813 net08208 net08202 vdd vdd nmos L=40e-9 W=180e-9
m1812 net08208 net08201 vdd vdd nmos L=40e-9 W=180e-9
m1811 net08239 net08232 vdd vdd nmos L=40e-9 W=180e-9
m1810 net08082 net08076 vdd vdd nmos L=40e-9 W=180e-9
m1809 net08082 net08075 vdd vdd nmos L=40e-9 W=180e-9
m1808 net08520 net08513 vdd vdd nmos L=40e-9 W=180e-9
m1807 net08520 net08514 vdd vdd nmos L=40e-9 W=180e-9
m1806 net08365 net08358 vdd vdd nmos L=40e-9 W=180e-9
m1805 net08365 net08359 vdd vdd nmos L=40e-9 W=180e-9
m1804 net08396 net08389 vdd vdd nmos L=40e-9 W=180e-9
m1803 net08396 net08390 vdd vdd nmos L=40e-9 W=180e-9
m1802 net08427 net08420 vdd vdd nmos L=40e-9 W=180e-9
m1801 net08427 net08421 vdd vdd nmos L=40e-9 W=180e-9
m1800 net08458 net08451 vdd vdd nmos L=40e-9 W=180e-9
m1799 net08458 net08452 vdd vdd nmos L=40e-9 W=180e-9
m1798 net08489 net08482 vdd vdd nmos L=40e-9 W=180e-9
m1797 net08489 net08483 vdd vdd nmos L=40e-9 W=180e-9
m1796 net08263 c48 vdd vdd nmos L=40e-9 W=180e-9
m1795 net08294 net08868 vdd vdd nmos L=40e-9 W=180e-9
m1794 net08325 c49 vdd vdd nmos L=40e-9 W=180e-9
m1793 net08108 c43 vdd vdd nmos L=40e-9 W=180e-9
m1792 net08139 c44 vdd vdd nmos L=40e-9 W=180e-9
m1791 net08170 c45 vdd vdd nmos L=40e-9 W=180e-9
m1790 net08201 c46 vdd vdd nmos L=40e-9 W=180e-9
m1789 net08232 c47 vdd vdd nmos L=40e-9 W=180e-9
m1788 net08075 c42 vdd vdd nmos L=40e-9 W=180e-9
m1787 net08513 c55 vdd vdd nmos L=40e-9 W=180e-9
m1786 net08358 c50 vdd vdd nmos L=40e-9 W=180e-9
m1785 net08389 c51 vdd vdd nmos L=40e-9 W=180e-9
m1784 net08420 c52 vdd vdd nmos L=40e-9 W=180e-9
m1783 net08451 c53 vdd vdd nmos L=40e-9 W=180e-9
m1782 net08482 c54 vdd vdd nmos L=40e-9 W=180e-9
m1743 net08359 net08334 vdd vdd nmos L=40e-9 W=180e-9
m1742 net08295 net08270 vdd vdd nmos L=40e-9 W=180e-9
m1741 net08295 net08272 vdd vdd nmos L=40e-9 W=180e-9
m1740 net08326 net08303 vdd vdd nmos L=40e-9 W=180e-9
m1739 net08326 net08301 vdd vdd nmos L=40e-9 W=180e-9
m1738 net08359 net08332 vdd vdd nmos L=40e-9 W=180e-9
m1736 net08140 net08117 vdd vdd nmos L=40e-9 W=180e-9
m1735 net08140 net08115 vdd vdd nmos L=40e-9 W=180e-9
m1734 net08171 net08148 vdd vdd nmos L=40e-9 W=180e-9
m1733 net08171 net08146 vdd vdd nmos L=40e-9 W=180e-9
m1732 net08202 net08177 vdd vdd nmos L=40e-9 W=180e-9
m1731 net08202 net08179 vdd vdd nmos L=40e-9 W=180e-9
m1730 net08233 net08210 vdd vdd nmos L=40e-9 W=180e-9
m1729 net08233 net08208 vdd vdd nmos L=40e-9 W=180e-9
m1728 net08264 net08239 vdd vdd nmos L=40e-9 W=180e-9
m1727 net08264 net08241 vdd vdd nmos L=40e-9 W=180e-9
m1726 net08109 net08084 vdd vdd nmos L=40e-9 W=180e-9
m1725 net08109 net08082 vdd vdd nmos L=40e-9 W=180e-9
m1718 net08545 net08520 vdd vdd nmos L=40e-9 W=180e-9
m1717 net08545 net08522 vdd vdd nmos L=40e-9 W=180e-9
m1716 net08390 net08365 vdd vdd nmos L=40e-9 W=180e-9
m1715 net08390 net08367 vdd vdd nmos L=40e-9 W=180e-9
m1714 net08421 net08396 vdd vdd nmos L=40e-9 W=180e-9
m1713 net08421 net08398 vdd vdd nmos L=40e-9 W=180e-9
m1712 net08452 net08427 vdd vdd nmos L=40e-9 W=180e-9
m1711 net08452 net08429 vdd vdd nmos L=40e-9 W=180e-9
m1710 net08483 net08458 vdd vdd nmos L=40e-9 W=180e-9
m1709 net08483 net08460 vdd vdd nmos L=40e-9 W=180e-9
m1708 net08514 net08489 vdd vdd nmos L=40e-9 W=180e-9
m1707 net08514 net08491 vdd vdd nmos L=40e-9 W=180e-9
m1688 net07832 net07825 vdd vdd nmos L=40e-9 W=180e-9
m1687 net07801 net07794 vdd vdd nmos L=40e-9 W=180e-9
m1686 net07801 net07795 vdd vdd nmos L=40e-9 W=180e-9
m1685 net07832 net07826 vdd vdd nmos L=40e-9 W=180e-9
m1684 net07770 net07764 vdd vdd nmos L=40e-9 W=180e-9
m1683 net07770 net07763 vdd vdd nmos L=40e-9 W=180e-9
m1682 net07739 net07732 vdd vdd nmos L=40e-9 W=180e-9
m1681 net07708 net07701 vdd vdd nmos L=40e-9 W=180e-9
m1680 net07708 net07702 vdd vdd nmos L=40e-9 W=180e-9
m1679 net07739 net07733 vdd vdd nmos L=40e-9 W=180e-9
m1678 net07677 net07671 vdd vdd nmos L=40e-9 W=180e-9
m1677 net07677 net07670 vdd vdd nmos L=40e-9 W=180e-9
m1676 net07646 net07639 vdd vdd nmos L=40e-9 W=180e-9
m1675 net07646 net07640 vdd vdd nmos L=40e-9 W=180e-9
m1674 net07615 net07608 vdd vdd nmos L=40e-9 W=180e-9
m1673 net07615 net07609 vdd vdd nmos L=40e-9 W=180e-9
m1672 net08051 net08045 vdd vdd nmos L=40e-9 W=180e-9
m1671 net08051 net08044 vdd vdd nmos L=40e-9 W=180e-9
m1670 net08020 net08014 vdd vdd nmos L=40e-9 W=180e-9
m1669 net08020 net08013 vdd vdd nmos L=40e-9 W=180e-9
m1668 net07989 net07983 vdd vdd nmos L=40e-9 W=180e-9
m1667 net07989 net07982 vdd vdd nmos L=40e-9 W=180e-9
m1666 net07958 net07952 vdd vdd nmos L=40e-9 W=180e-9
m1665 net07958 net07951 vdd vdd nmos L=40e-9 W=180e-9
m1664 net07927 net07921 vdd vdd nmos L=40e-9 W=180e-9
m1663 net07927 net07920 vdd vdd nmos L=40e-9 W=180e-9
m1662 net07896 net07890 vdd vdd nmos L=40e-9 W=180e-9
m1661 net07896 net07889 vdd vdd nmos L=40e-9 W=180e-9
m1660 net07865 net07859 vdd vdd nmos L=40e-9 W=180e-9
m1659 net07865 net07858 vdd vdd nmos L=40e-9 W=180e-9
m1658 net07825 c35 vdd vdd nmos L=40e-9 W=180e-9
m1657 net07794 c34 vdd vdd nmos L=40e-9 W=180e-9
m1656 net07763 c33 vdd vdd nmos L=40e-9 W=180e-9
m1655 net07732 net08836 vdd vdd nmos L=40e-9 W=180e-9
m1654 net07701 c32 vdd vdd nmos L=40e-9 W=180e-9
m1653 net07670 c31 vdd vdd nmos L=40e-9 W=180e-9
m1652 net07639 c30 vdd vdd nmos L=40e-9 W=180e-9
m1651 net07608 c29 vdd vdd nmos L=40e-9 W=180e-9
m1650 net08044 c41 vdd vdd nmos L=40e-9 W=180e-9
m1649 net08013 net08852 vdd vdd nmos L=40e-9 W=180e-9
m1648 net07982 c40 vdd vdd nmos L=40e-9 W=180e-9
m1647 net07951 c39 vdd vdd nmos L=40e-9 W=180e-9
m1646 net07920 c38 vdd vdd nmos L=40e-9 W=180e-9
m1645 net07889 c37 vdd vdd nmos L=40e-9 W=180e-9
m1644 net07858 c36 vdd vdd nmos L=40e-9 W=180e-9
m1610 net07859 net07832 vdd vdd nmos L=40e-9 W=180e-9
m1609 net07826 net07801 vdd vdd nmos L=40e-9 W=180e-9
m1608 net07826 net07803 vdd vdd nmos L=40e-9 W=180e-9
m1607 net07795 net07772 vdd vdd nmos L=40e-9 W=180e-9
m1606 net07795 net07770 vdd vdd nmos L=40e-9 W=180e-9
m1605 net07859 net07834 vdd vdd nmos L=40e-9 W=180e-9
m1599 net07764 net07741 vdd vdd nmos L=40e-9 W=180e-9
m1598 net07764 net07739 vdd vdd nmos L=40e-9 W=180e-9
m1597 net07733 net07708 vdd vdd nmos L=40e-9 W=180e-9
m1596 net07733 net07710 vdd vdd nmos L=40e-9 W=180e-9
m1595 net07702 net07679 vdd vdd nmos L=40e-9 W=180e-9
m1594 net07702 net07677 vdd vdd nmos L=40e-9 W=180e-9
m1593 net07671 net07646 vdd vdd nmos L=40e-9 W=180e-9
m1592 net07671 net07648 vdd vdd nmos L=40e-9 W=180e-9
m1591 net07640 net07615 vdd vdd nmos L=40e-9 W=180e-9
m1590 net07640 net07617 vdd vdd nmos L=40e-9 W=180e-9
m1587 net08076 net08053 vdd vdd nmos L=40e-9 W=180e-9
m1586 net08076 net08051 vdd vdd nmos L=40e-9 W=180e-9
m1585 net08045 net08022 vdd vdd nmos L=40e-9 W=180e-9
m1584 net08045 net08020 vdd vdd nmos L=40e-9 W=180e-9
m1578 net08014 net07991 vdd vdd nmos L=40e-9 W=180e-9
m1577 net08014 net07989 vdd vdd nmos L=40e-9 W=180e-9
m1576 net07983 net07960 vdd vdd nmos L=40e-9 W=180e-9
m1575 net07983 net07958 vdd vdd nmos L=40e-9 W=180e-9
m1574 net07952 net07929 vdd vdd nmos L=40e-9 W=180e-9
m1573 net07952 net07927 vdd vdd nmos L=40e-9 W=180e-9
m1572 net07921 net07898 vdd vdd nmos L=40e-9 W=180e-9
m1571 net07921 net07896 vdd vdd nmos L=40e-9 W=180e-9
m1570 net07890 net07867 vdd vdd nmos L=40e-9 W=180e-9
m1569 net07890 net07865 vdd vdd nmos L=40e-9 W=180e-9
m1543 net08553 c56 vdd vdd nmos L=40e-9 W=180e-9
m1542 net08553 net08528 vdd vdd nmos L=40e-9 W=180e-9
m1541 net08584 net08884 vdd vdd nmos L=40e-9 W=180e-9
m1540 net08584 net08559 vdd vdd nmos L=40e-9 W=180e-9
m1535 net08547 net08541 vdd vdd nmos L=40e-9 W=180e-9
m1534 net08547 net08528 vdd vdd nmos L=40e-9 W=180e-9
m1533 net08578 net08559 vdd vdd nmos L=40e-9 W=180e-9
m1532 net08578 net08572 vdd vdd nmos L=40e-9 W=180e-9
m1531 net08572 net08884 vdd vdd nmos L=40e-9 W=180e-9
m1530 net08541 c56 vdd vdd nmos L=40e-9 W=180e-9
m1523 net08559 net08549 vdd vdd nmos L=40e-9 W=180e-9
m1522 net08593 net08580 vdd vdd nmos L=40e-9 W=180e-9
m1521 net08593 net08578 vdd vdd nmos L=40e-9 W=180e-9
m1520 net08559 net08547 vdd vdd nmos L=40e-9 W=180e-9
m1513 net08272 c48 vdd vdd nmos L=40e-9 W=180e-9
m1512 net08272 net08247 vdd vdd nmos L=40e-9 W=180e-9
m1511 net08303 net08278 vdd vdd nmos L=40e-9 W=180e-9
m1510 net08303 net08868 vdd vdd nmos L=40e-9 W=180e-9
m1509 net08334 c49 vdd vdd nmos L=40e-9 W=180e-9
m1508 net08334 net08309 vdd vdd nmos L=40e-9 W=180e-9
m1506 net08117 net08093 vdd vdd nmos L=40e-9 W=180e-9
m1505 net08117 c43 vdd vdd nmos L=40e-9 W=180e-9
m1504 net08148 net08123 vdd vdd nmos L=40e-9 W=180e-9
m1503 net08148 c44 vdd vdd nmos L=40e-9 W=180e-9
m1502 net08179 c45 vdd vdd nmos L=40e-9 W=180e-9
m1501 net08179 net08154 vdd vdd nmos L=40e-9 W=180e-9
m1500 net08210 net08185 vdd vdd nmos L=40e-9 W=180e-9
m1499 net08210 c46 vdd vdd nmos L=40e-9 W=180e-9
m1498 net08241 c47 vdd vdd nmos L=40e-9 W=180e-9
m1497 net08241 net08216 vdd vdd nmos L=40e-9 W=180e-9
m1491 net08084 net08059 vdd vdd nmos L=40e-9 W=180e-9
m1490 net08084 c42 vdd vdd nmos L=40e-9 W=180e-9
m1489 net08522 c55 vdd vdd nmos L=40e-9 W=180e-9
m1488 net08522 net08497 vdd vdd nmos L=40e-9 W=180e-9
m1487 net08367 c50 vdd vdd nmos L=40e-9 W=180e-9
m1486 net08367 net08343 vdd vdd nmos L=40e-9 W=180e-9
m1485 net08398 c51 vdd vdd nmos L=40e-9 W=180e-9
m1484 net08398 net08373 vdd vdd nmos L=40e-9 W=180e-9
m1483 net08429 c52 vdd vdd nmos L=40e-9 W=180e-9
m1482 net08429 net08404 vdd vdd nmos L=40e-9 W=180e-9
m1481 net08460 c53 vdd vdd nmos L=40e-9 W=180e-9
m1480 net08460 net08435 vdd vdd nmos L=40e-9 W=180e-9
m1479 net08491 c54 vdd vdd nmos L=40e-9 W=180e-9
m1478 net08491 net08466 vdd vdd nmos L=40e-9 W=180e-9
m1447 net08266 net08260 vdd vdd nmos L=40e-9 W=180e-9
m1446 net08266 net08247 vdd vdd nmos L=40e-9 W=180e-9
m1445 net08297 net08278 vdd vdd nmos L=40e-9 W=180e-9
m1444 net08297 net08291 vdd vdd nmos L=40e-9 W=180e-9
m1443 net08328 net08322 vdd vdd nmos L=40e-9 W=180e-9
m1442 net08328 net08309 vdd vdd nmos L=40e-9 W=180e-9
m1441 net08111 net08093 vdd vdd nmos L=40e-9 W=180e-9
m1440 net08111 net08105 vdd vdd nmos L=40e-9 W=180e-9
m1439 net08142 net08123 vdd vdd nmos L=40e-9 W=180e-9
m1438 net08142 net08136 vdd vdd nmos L=40e-9 W=180e-9
m1437 net08173 net08167 vdd vdd nmos L=40e-9 W=180e-9
m1436 net08173 net08154 vdd vdd nmos L=40e-9 W=180e-9
m1435 net08204 net08185 vdd vdd nmos L=40e-9 W=180e-9
m1434 net08204 net08198 vdd vdd nmos L=40e-9 W=180e-9
m1433 net08235 net08229 vdd vdd nmos L=40e-9 W=180e-9
m1432 net08235 net08216 vdd vdd nmos L=40e-9 W=180e-9
m1431 net08078 net08072 vdd vdd nmos L=40e-9 W=180e-9
m1430 net08078 net08059 vdd vdd nmos L=40e-9 W=180e-9
m1429 net08516 net08497 vdd vdd nmos L=40e-9 W=180e-9
m1428 net08516 net08510 vdd vdd nmos L=40e-9 W=180e-9
m1427 net08485 net08466 vdd vdd nmos L=40e-9 W=180e-9
m1426 net08485 net08479 vdd vdd nmos L=40e-9 W=180e-9
m1425 net08454 net08448 vdd vdd nmos L=40e-9 W=180e-9
m1424 net08454 net08435 vdd vdd nmos L=40e-9 W=180e-9
m1423 net08423 net08404 vdd vdd nmos L=40e-9 W=180e-9
m1422 net08423 net08417 vdd vdd nmos L=40e-9 W=180e-9
m1421 net08392 net08386 vdd vdd nmos L=40e-9 W=180e-9
m1420 net08392 net08373 vdd vdd nmos L=40e-9 W=180e-9
m1419 net08361 net08355 vdd vdd nmos L=40e-9 W=180e-9
m1418 net08361 net08343 vdd vdd nmos L=40e-9 W=180e-9
m1417 net08260 c48 vdd vdd nmos L=40e-9 W=180e-9
m1416 net08291 net08868 vdd vdd nmos L=40e-9 W=180e-9
m1415 net08322 c49 vdd vdd nmos L=40e-9 W=180e-9
m1414 net08105 c43 vdd vdd nmos L=40e-9 W=180e-9
m1413 net08136 c44 vdd vdd nmos L=40e-9 W=180e-9
m1412 net08167 c45 vdd vdd nmos L=40e-9 W=180e-9
m1411 net08198 c46 vdd vdd nmos L=40e-9 W=180e-9
m1410 net08229 c47 vdd vdd nmos L=40e-9 W=180e-9
m1409 net08072 c42 vdd vdd nmos L=40e-9 W=180e-9
m1408 net08510 c55 vdd vdd nmos L=40e-9 W=180e-9
m1407 net08479 c54 vdd vdd nmos L=40e-9 W=180e-9
m1406 net08448 c53 vdd vdd nmos L=40e-9 W=180e-9
m1405 net08417 c52 vdd vdd nmos L=40e-9 W=180e-9
m1404 net08386 c51 vdd vdd nmos L=40e-9 W=180e-9
m1403 net08355 c50 vdd vdd nmos L=40e-9 W=180e-9
m1364 net08278 net08266 vdd vdd nmos L=40e-9 W=180e-9
m1363 net08278 net08268 vdd vdd nmos L=40e-9 W=180e-9
m1362 net08309 net08299 vdd vdd nmos L=40e-9 W=180e-9
m1361 net08309 net08297 vdd vdd nmos L=40e-9 W=180e-9
m1360 net08343 net08328 vdd vdd nmos L=40e-9 W=180e-9
m1359 net08343 net08330 vdd vdd nmos L=40e-9 W=180e-9
m1357 net08123 net08111 vdd vdd nmos L=40e-9 W=180e-9
m1356 net08154 net08144 vdd vdd nmos L=40e-9 W=180e-9
m1355 net08154 net08142 vdd vdd nmos L=40e-9 W=180e-9
m1354 net08185 net08173 vdd vdd nmos L=40e-9 W=180e-9
m1353 net08185 net08175 vdd vdd nmos L=40e-9 W=180e-9
m1352 net08216 net08206 vdd vdd nmos L=40e-9 W=180e-9
m1351 net08216 net08204 vdd vdd nmos L=40e-9 W=180e-9
m1350 net08247 net08235 vdd vdd nmos L=40e-9 W=180e-9
m1349 net08247 net08237 vdd vdd nmos L=40e-9 W=180e-9
m1348 net08123 net08113 vdd vdd nmos L=40e-9 W=180e-9
m1347 net08093 net08078 vdd vdd nmos L=40e-9 W=180e-9
m1346 net08093 net08080 vdd vdd nmos L=40e-9 W=180e-9
m1344 net08528 net08518 vdd vdd nmos L=40e-9 W=180e-9
m1343 net08528 net08516 vdd vdd nmos L=40e-9 W=180e-9
m1337 net08497 net08487 vdd vdd nmos L=40e-9 W=180e-9
m1336 net08497 net08485 vdd vdd nmos L=40e-9 W=180e-9
m1335 net08466 net08454 vdd vdd nmos L=40e-9 W=180e-9
m1334 net08466 net08456 vdd vdd nmos L=40e-9 W=180e-9
m1333 net08435 net08425 vdd vdd nmos L=40e-9 W=180e-9
m1332 net08435 net08423 vdd vdd nmos L=40e-9 W=180e-9
m1331 net08404 net08392 vdd vdd nmos L=40e-9 W=180e-9
m1330 net08404 net08394 vdd vdd nmos L=40e-9 W=180e-9
m1329 net08373 net08361 vdd vdd nmos L=40e-9 W=180e-9
m1328 net08373 net08363 vdd vdd nmos L=40e-9 W=180e-9
m1325 net07834 net07809 vdd vdd nmos L=40e-9 W=180e-9
m1324 net07834 c35 vdd vdd nmos L=40e-9 W=180e-9
m1323 net07803 c34 vdd vdd nmos L=40e-9 W=180e-9
m1322 net07803 net07778 vdd vdd nmos L=40e-9 W=180e-9
m1321 net07772 net07747 vdd vdd nmos L=40e-9 W=180e-9
m1320 net07772 c33 vdd vdd nmos L=40e-9 W=180e-9
m1314 net07741 net07716 vdd vdd nmos L=40e-9 W=180e-9
m1313 net07741 net08836 vdd vdd nmos L=40e-9 W=180e-9
m1312 net07710 c32 vdd vdd nmos L=40e-9 W=180e-9
m1311 net07710 net07685 vdd vdd nmos L=40e-9 W=180e-9
m1310 net07679 net07654 vdd vdd nmos L=40e-9 W=180e-9
m1309 net07679 c31 vdd vdd nmos L=40e-9 W=180e-9
m1308 net07648 c30 vdd vdd nmos L=40e-9 W=180e-9
m1307 net07648 net07623 vdd vdd nmos L=40e-9 W=180e-9
m1306 net07617 c29 vdd vdd nmos L=40e-9 W=180e-9
m1305 net07617 net07593 vdd vdd nmos L=40e-9 W=180e-9
m1304 net08053 net08028 vdd vdd nmos L=40e-9 W=180e-9
m1303 net08053 c41 vdd vdd nmos L=40e-9 W=180e-9
m1302 net08022 net07997 vdd vdd nmos L=40e-9 W=180e-9
m1301 net08022 net08852 vdd vdd nmos L=40e-9 W=180e-9
m1300 net07991 net07966 vdd vdd nmos L=40e-9 W=180e-9
m1299 net07991 c40 vdd vdd nmos L=40e-9 W=180e-9
m1298 net07960 net07935 vdd vdd nmos L=40e-9 W=180e-9
m1297 net07960 c39 vdd vdd nmos L=40e-9 W=180e-9
m1296 net07929 net07904 vdd vdd nmos L=40e-9 W=180e-9
m1295 net07929 c38 vdd vdd nmos L=40e-9 W=180e-9
m1294 net07898 net07873 vdd vdd nmos L=40e-9 W=180e-9
m1293 net07898 c37 vdd vdd nmos L=40e-9 W=180e-9
m1292 net07867 net07843 vdd vdd nmos L=40e-9 W=180e-9
m1291 net07867 c36 vdd vdd nmos L=40e-9 W=180e-9
m1260 net07828 net07809 vdd vdd nmos L=40e-9 W=180e-9
m1259 net07828 net07822 vdd vdd nmos L=40e-9 W=180e-9
m1258 net07797 net07791 vdd vdd nmos L=40e-9 W=180e-9
m1257 net07797 net07778 vdd vdd nmos L=40e-9 W=180e-9
m1256 net07766 net07747 vdd vdd nmos L=40e-9 W=180e-9
m1255 net07766 net07760 vdd vdd nmos L=40e-9 W=180e-9
m1254 net07735 net07716 vdd vdd nmos L=40e-9 W=180e-9
m1253 net07735 net07729 vdd vdd nmos L=40e-9 W=180e-9
m1252 net07704 net07698 vdd vdd nmos L=40e-9 W=180e-9
m1251 net07704 net07685 vdd vdd nmos L=40e-9 W=180e-9
m1250 net07673 net07654 vdd vdd nmos L=40e-9 W=180e-9
m1249 net07673 net07667 vdd vdd nmos L=40e-9 W=180e-9
m1248 net07642 net07636 vdd vdd nmos L=40e-9 W=180e-9
m1247 net07642 net07623 vdd vdd nmos L=40e-9 W=180e-9
m1246 net07611 net07605 vdd vdd nmos L=40e-9 W=180e-9
m1245 net07611 net07593 vdd vdd nmos L=40e-9 W=180e-9
m1244 net08016 net08010 vdd vdd nmos L=40e-9 W=180e-9
m1243 net08016 net07997 vdd vdd nmos L=40e-9 W=180e-9
m1242 net08047 net08028 vdd vdd nmos L=40e-9 W=180e-9
m1241 net08047 net08041 vdd vdd nmos L=40e-9 W=180e-9
m1240 net07861 net07843 vdd vdd nmos L=40e-9 W=180e-9
m1239 net07861 net07855 vdd vdd nmos L=40e-9 W=180e-9
m1238 net07892 net07873 vdd vdd nmos L=40e-9 W=180e-9
m1237 net07892 net07886 vdd vdd nmos L=40e-9 W=180e-9
m1236 net07923 net07917 vdd vdd nmos L=40e-9 W=180e-9
m1235 net07923 net07904 vdd vdd nmos L=40e-9 W=180e-9
m1234 net07954 net07935 vdd vdd nmos L=40e-9 W=180e-9
m1233 net07954 net07948 vdd vdd nmos L=40e-9 W=180e-9
m1232 net07985 net07979 vdd vdd nmos L=40e-9 W=180e-9
m1231 net07985 net07966 vdd vdd nmos L=40e-9 W=180e-9
m1230 net07822 c35 vdd vdd nmos L=40e-9 W=180e-9
m1229 net07791 c34 vdd vdd nmos L=40e-9 W=180e-9
m1228 net07760 c33 vdd vdd nmos L=40e-9 W=180e-9
m1227 net07729 net08836 vdd vdd nmos L=40e-9 W=180e-9
m1226 net07698 c32 vdd vdd nmos L=40e-9 W=180e-9
m1225 net07667 c31 vdd vdd nmos L=40e-9 W=180e-9
m1224 net07636 c30 vdd vdd nmos L=40e-9 W=180e-9
m1223 net07605 c29 vdd vdd nmos L=40e-9 W=180e-9
m1222 net08010 net08852 vdd vdd nmos L=40e-9 W=180e-9
m1221 net08041 c41 vdd vdd nmos L=40e-9 W=180e-9
m1220 net07855 c36 vdd vdd nmos L=40e-9 W=180e-9
m1219 net07886 c37 vdd vdd nmos L=40e-9 W=180e-9
m1218 net07917 c38 vdd vdd nmos L=40e-9 W=180e-9
m1217 net07948 c39 vdd vdd nmos L=40e-9 W=180e-9
m1216 net07979 c40 vdd vdd nmos L=40e-9 W=180e-9
m1182 net07843 net07830 vdd vdd nmos L=40e-9 W=180e-9
m1181 net07843 net07828 vdd vdd nmos L=40e-9 W=180e-9
m1180 net07809 net07797 vdd vdd nmos L=40e-9 W=180e-9
m1179 net07809 net07799 vdd vdd nmos L=40e-9 W=180e-9
m1178 net07778 net07768 vdd vdd nmos L=40e-9 W=180e-9
m1177 net07778 net07766 vdd vdd nmos L=40e-9 W=180e-9
m1171 net07747 net07737 vdd vdd nmos L=40e-9 W=180e-9
m1170 net07747 net07735 vdd vdd nmos L=40e-9 W=180e-9
m1169 net07716 net07704 vdd vdd nmos L=40e-9 W=180e-9
m1168 net07716 net07706 vdd vdd nmos L=40e-9 W=180e-9
m1167 net07685 net07675 vdd vdd nmos L=40e-9 W=180e-9
m1166 net07685 net07673 vdd vdd nmos L=40e-9 W=180e-9
m1165 net07654 net07642 vdd vdd nmos L=40e-9 W=180e-9
m1164 net07654 net07644 vdd vdd nmos L=40e-9 W=180e-9
m1163 net07623 net07611 vdd vdd nmos L=40e-9 W=180e-9
m1162 net07623 net07613 vdd vdd nmos L=40e-9 W=180e-9
m1154 net08028 net08016 vdd vdd nmos L=40e-9 W=180e-9
m1153 net08028 net08018 vdd vdd nmos L=40e-9 W=180e-9
m1152 net08059 net08049 vdd vdd nmos L=40e-9 W=180e-9
m1151 net08059 net08047 vdd vdd nmos L=40e-9 W=180e-9
m1150 net07873 net07863 vdd vdd nmos L=40e-9 W=180e-9
m1149 net07873 net07861 vdd vdd nmos L=40e-9 W=180e-9
m1148 net07904 net07894 vdd vdd nmos L=40e-9 W=180e-9
m1147 net07904 net07892 vdd vdd nmos L=40e-9 W=180e-9
m1146 net07935 net07923 vdd vdd nmos L=40e-9 W=180e-9
m1145 net07935 net07925 vdd vdd nmos L=40e-9 W=180e-9
m1144 net07966 net07956 vdd vdd nmos L=40e-9 W=180e-9
m1143 net07966 net07954 vdd vdd nmos L=40e-9 W=180e-9
m1142 net07997 net07985 vdd vdd nmos L=40e-9 W=180e-9
m1141 net07997 net07987 vdd vdd nmos L=40e-9 W=180e-9
m1136 net08549 c56 vdd vdd nmos L=40e-9 W=180e-9
m1135 net08549 net08545 vdd vdd nmos L=40e-9 W=180e-9
m1134 net08580 net08576 vdd vdd nmos L=40e-9 W=180e-9
m1133 net08580 net08884 vdd vdd nmos L=40e-9 W=180e-9
m1104 net08268 c48 vdd vdd nmos L=40e-9 W=180e-9
m1103 net08268 net08264 vdd vdd nmos L=40e-9 W=180e-9
m1102 net08299 net08295 vdd vdd nmos L=40e-9 W=180e-9
m1101 net08299 net08868 vdd vdd nmos L=40e-9 W=180e-9
m1100 net08330 c49 vdd vdd nmos L=40e-9 W=180e-9
m1099 net08330 net08326 vdd vdd nmos L=40e-9 W=180e-9
m1097 net08113 net08109 vdd vdd nmos L=40e-9 W=180e-9
m1096 net08113 c43 vdd vdd nmos L=40e-9 W=180e-9
m1095 net08144 net08140 vdd vdd nmos L=40e-9 W=180e-9
m1094 net08144 c44 vdd vdd nmos L=40e-9 W=180e-9
m1093 net08175 c45 vdd vdd nmos L=40e-9 W=180e-9
m1092 net08175 net08171 vdd vdd nmos L=40e-9 W=180e-9
m1091 net08206 net08202 vdd vdd nmos L=40e-9 W=180e-9
m1090 net08206 c46 vdd vdd nmos L=40e-9 W=180e-9
m1089 net08237 c47 vdd vdd nmos L=40e-9 W=180e-9
m1088 net08237 net08233 vdd vdd nmos L=40e-9 W=180e-9
m1082 net08080 c42 vdd vdd nmos L=40e-9 W=180e-9
m1081 net08080 net08076 vdd vdd nmos L=40e-9 W=180e-9
m1080 net08518 net08514 vdd vdd nmos L=40e-9 W=180e-9
m1079 net08518 c55 vdd vdd nmos L=40e-9 W=180e-9
m1078 net08487 net08483 vdd vdd nmos L=40e-9 W=180e-9
m1077 net08487 c54 vdd vdd nmos L=40e-9 W=180e-9
m1076 net08456 c53 vdd vdd nmos L=40e-9 W=180e-9
m1075 net08456 net08452 vdd vdd nmos L=40e-9 W=180e-9
m1074 net08425 net08421 vdd vdd nmos L=40e-9 W=180e-9
m1073 net08425 c52 vdd vdd nmos L=40e-9 W=180e-9
m1072 net08394 c51 vdd vdd nmos L=40e-9 W=180e-9
m1071 net08394 net08390 vdd vdd nmos L=40e-9 W=180e-9
m1070 net08363 c50 vdd vdd nmos L=40e-9 W=180e-9
m1069 net08363 net08359 vdd vdd nmos L=40e-9 W=180e-9
m1013 net07830 net07826 vdd vdd nmos L=40e-9 W=180e-9
m1012 net07830 c35 vdd vdd nmos L=40e-9 W=180e-9
m1011 net07799 c34 vdd vdd nmos L=40e-9 W=180e-9
m1010 net07799 net07795 vdd vdd nmos L=40e-9 W=180e-9
m1009 net07768 net07764 vdd vdd nmos L=40e-9 W=180e-9
m1008 net07768 c33 vdd vdd nmos L=40e-9 W=180e-9
m1002 net07737 net07733 vdd vdd nmos L=40e-9 W=180e-9
m1001 net07737 net08836 vdd vdd nmos L=40e-9 W=180e-9
m1000 net07706 c32 vdd vdd nmos L=40e-9 W=180e-9
m999 net07706 net07702 vdd vdd nmos L=40e-9 W=180e-9
m998 net07675 net07671 vdd vdd nmos L=40e-9 W=180e-9
m997 net07675 c31 vdd vdd nmos L=40e-9 W=180e-9
m996 net07644 c30 vdd vdd nmos L=40e-9 W=180e-9
m995 net07644 net07640 vdd vdd nmos L=40e-9 W=180e-9
m994 net07613 c29 vdd vdd nmos L=40e-9 W=180e-9
m993 net07613 net07609 vdd vdd nmos L=40e-9 W=180e-9
m992 net08018 net08852 vdd vdd nmos L=40e-9 W=180e-9
m991 net08018 net08014 vdd vdd nmos L=40e-9 W=180e-9
m990 net08049 net08045 vdd vdd nmos L=40e-9 W=180e-9
m989 net08049 c41 vdd vdd nmos L=40e-9 W=180e-9
m988 net07863 net07859 vdd vdd nmos L=40e-9 W=180e-9
m987 net07863 c36 vdd vdd nmos L=40e-9 W=180e-9
m986 net07894 net07890 vdd vdd nmos L=40e-9 W=180e-9
m985 net07894 c37 vdd vdd nmos L=40e-9 W=180e-9
m984 net07925 c38 vdd vdd nmos L=40e-9 W=180e-9
m983 net07925 net07921 vdd vdd nmos L=40e-9 W=180e-9
m982 net07956 net07952 vdd vdd nmos L=40e-9 W=180e-9
m981 net07956 c39 vdd vdd nmos L=40e-9 W=180e-9
m980 net07987 c40 vdd vdd nmos L=40e-9 W=180e-9
m979 net07987 net07983 vdd vdd nmos L=40e-9 W=180e-9
m948 net07609 net07584 vdd vdd nmos L=40e-9 W=180e-9
m945 net07609 net07582 vdd vdd nmos L=40e-9 W=180e-9
m944 net07584 net07559 vdd vdd nmos L=40e-9 W=180e-9
m943 net07582 net07576 vdd vdd nmos L=40e-9 W=180e-9
m938 net07584 c28 vdd vdd nmos L=40e-9 W=180e-9
m937 net07582 net07575 vdd vdd nmos L=40e-9 W=180e-9
m935 net07575 c28 vdd vdd nmos L=40e-9 W=180e-9
m934 net07576 net07552 vdd vdd nmos L=40e-9 W=180e-9
m931 net07576 net07550 vdd vdd nmos L=40e-9 W=180e-9
m930 net07552 net07527 vdd vdd nmos L=40e-9 W=180e-9
m929 net07550 net07544 vdd vdd nmos L=40e-9 W=180e-9
m924 net07552 c27 vdd vdd nmos L=40e-9 W=180e-9
m923 net07550 net07543 vdd vdd nmos L=40e-9 W=180e-9
m921 net07543 c27 vdd vdd nmos L=40e-9 W=180e-9
m920 net07544 net07520 vdd vdd nmos L=40e-9 W=180e-9
m917 net07544 net07518 vdd vdd nmos L=40e-9 W=180e-9
m916 net07520 net07494 vdd vdd nmos L=40e-9 W=180e-9
m915 net07518 net07511 vdd vdd nmos L=40e-9 W=180e-9
m910 net07520 c26 vdd vdd nmos L=40e-9 W=180e-9
m909 net07518 net07510 vdd vdd nmos L=40e-9 W=180e-9
m907 net07510 c26 vdd vdd nmos L=40e-9 W=180e-9
m906 net07511 net07488 vdd vdd nmos L=40e-9 W=180e-9
m903 net07511 net07486 vdd vdd nmos L=40e-9 W=180e-9
m902 net07488 net07463 vdd vdd nmos L=40e-9 W=180e-9
m901 net07486 net07480 vdd vdd nmos L=40e-9 W=180e-9
m896 net07488 c25 vdd vdd nmos L=40e-9 W=180e-9
m895 net07486 net07479 vdd vdd nmos L=40e-9 W=180e-9
m893 net07479 c25 vdd vdd nmos L=40e-9 W=180e-9
m892 net07480 net07457 vdd vdd nmos L=40e-9 W=180e-9
m889 net07480 net07455 vdd vdd nmos L=40e-9 W=180e-9
m888 net07457 net07432 vdd vdd nmos L=40e-9 W=180e-9
m887 net07455 net07449 vdd vdd nmos L=40e-9 W=180e-9
m882 net07457 net08819 vdd vdd nmos L=40e-9 W=180e-9
m881 net07455 net07448 vdd vdd nmos L=40e-9 W=180e-9
m879 net07448 net08819 vdd vdd nmos L=40e-9 W=180e-9
m878 net07449 net07426 vdd vdd nmos L=40e-9 W=180e-9
m875 net07449 net07424 vdd vdd nmos L=40e-9 W=180e-9
m874 net07426 net07401 vdd vdd nmos L=40e-9 W=180e-9
m873 net07424 net07418 vdd vdd nmos L=40e-9 W=180e-9
m868 net07426 c24 vdd vdd nmos L=40e-9 W=180e-9
m867 net07424 net07417 vdd vdd nmos L=40e-9 W=180e-9
m865 net07417 c24 vdd vdd nmos L=40e-9 W=180e-9
m864 net07418 net07395 vdd vdd nmos L=40e-9 W=180e-9
m861 net07418 net07393 vdd vdd nmos L=40e-9 W=180e-9
m860 net07395 net07370 vdd vdd nmos L=40e-9 W=180e-9
m859 net07393 net07387 vdd vdd nmos L=40e-9 W=180e-9
m854 net07395 c23 vdd vdd nmos L=40e-9 W=180e-9
m853 net07393 net07386 vdd vdd nmos L=40e-9 W=180e-9
m851 net07386 c23 vdd vdd nmos L=40e-9 W=180e-9
m850 net07387 net07364 vdd vdd nmos L=40e-9 W=180e-9
m847 net07387 net07362 vdd vdd nmos L=40e-9 W=180e-9
m846 net07364 net07340 vdd vdd nmos L=40e-9 W=180e-9
m845 net07362 net07356 vdd vdd nmos L=40e-9 W=180e-9
m840 net07364 c22 vdd vdd nmos L=40e-9 W=180e-9
m839 net07362 net07355 vdd vdd nmos L=40e-9 W=180e-9
m837 net07355 c22 vdd vdd nmos L=40e-9 W=180e-9
m836 net07329 net07322 vdd vdd nmos L=40e-9 W=180e-9
m835 net07298 net07291 vdd vdd nmos L=40e-9 W=180e-9
m834 net07298 net07292 vdd vdd nmos L=40e-9 W=180e-9
m833 net07329 net07323 vdd vdd nmos L=40e-9 W=180e-9
m832 net07267 net07261 vdd vdd nmos L=40e-9 W=180e-9
m831 net07267 net07260 vdd vdd nmos L=40e-9 W=180e-9
m830 net07236 net07228 vdd vdd nmos L=40e-9 W=180e-9
m829 net07204 net07197 vdd vdd nmos L=40e-9 W=180e-9
m828 net07204 net07198 vdd vdd nmos L=40e-9 W=180e-9
m827 net07236 net07229 vdd vdd nmos L=40e-9 W=180e-9
m826 net07173 net07167 vdd vdd nmos L=40e-9 W=180e-9
m825 net07173 net07166 vdd vdd nmos L=40e-9 W=180e-9
m824 net07142 net07135 vdd vdd nmos L=40e-9 W=180e-9
m823 net07142 net07136 vdd vdd nmos L=40e-9 W=180e-9
m822 net07111 net07104 vdd vdd nmos L=40e-9 W=180e-9
m821 net07111 net07105 vdd vdd nmos L=40e-9 W=180e-9
m820 net07322 c21 vdd vdd nmos L=40e-9 W=180e-9
m819 net07291 c20 vdd vdd nmos L=40e-9 W=180e-9
m818 net07260 c19 vdd vdd nmos L=40e-9 W=180e-9
m817 net07228 c18 vdd vdd nmos L=40e-9 W=180e-9
m816 net07197 c17 vdd vdd nmos L=40e-9 W=180e-9
m815 net07166 net08803 vdd vdd nmos L=40e-9 W=180e-9
m814 net07135 c16 vdd vdd nmos L=40e-9 W=180e-9
m813 net07104 c15 vdd vdd nmos L=40e-9 W=180e-9
m793 net07356 net07329 vdd vdd nmos L=40e-9 W=180e-9
m792 net07323 net07298 vdd vdd nmos L=40e-9 W=180e-9
m791 net07323 net07300 vdd vdd nmos L=40e-9 W=180e-9
m790 net07292 net07269 vdd vdd nmos L=40e-9 W=180e-9
m789 net07292 net07267 vdd vdd nmos L=40e-9 W=180e-9
m788 net07356 net07331 vdd vdd nmos L=40e-9 W=180e-9
m782 net07261 net07238 vdd vdd nmos L=40e-9 W=180e-9
m781 net07261 net07236 vdd vdd nmos L=40e-9 W=180e-9
m780 net07229 net07204 vdd vdd nmos L=40e-9 W=180e-9
m779 net07229 net07206 vdd vdd nmos L=40e-9 W=180e-9
m778 net07198 net07175 vdd vdd nmos L=40e-9 W=180e-9
m777 net07198 net07173 vdd vdd nmos L=40e-9 W=180e-9
m776 net07167 net07142 vdd vdd nmos L=40e-9 W=180e-9
m775 net07167 net07144 vdd vdd nmos L=40e-9 W=180e-9
m774 net07136 net07111 vdd vdd nmos L=40e-9 W=180e-9
m773 net07136 net07113 vdd vdd nmos L=40e-9 W=180e-9
m756 net07331 net07306 vdd vdd nmos L=40e-9 W=180e-9
m755 net07331 c21 vdd vdd nmos L=40e-9 W=180e-9
m754 net07300 c20 vdd vdd nmos L=40e-9 W=180e-9
m753 net07300 net07275 vdd vdd nmos L=40e-9 W=180e-9
m752 net07269 net07244 vdd vdd nmos L=40e-9 W=180e-9
m751 net07269 c19 vdd vdd nmos L=40e-9 W=180e-9
m750 net07238 net07212 vdd vdd nmos L=40e-9 W=180e-9
m749 net07238 c18 vdd vdd nmos L=40e-9 W=180e-9
m748 net07206 c17 vdd vdd nmos L=40e-9 W=180e-9
m747 net07206 net07181 vdd vdd nmos L=40e-9 W=180e-9
m746 net07175 net07150 vdd vdd nmos L=40e-9 W=180e-9
m745 net07175 net08803 vdd vdd nmos L=40e-9 W=180e-9
m744 net07144 c16 vdd vdd nmos L=40e-9 W=180e-9
m743 net07144 net07119 vdd vdd nmos L=40e-9 W=180e-9
m742 net07113 c15 vdd vdd nmos L=40e-9 W=180e-9
m741 net07113 net07089 vdd vdd nmos L=40e-9 W=180e-9
m724 net07578 net07572 vdd vdd nmos L=40e-9 W=180e-9
m723 net07578 net07559 vdd vdd nmos L=40e-9 W=180e-9
m720 net07593 net07578 vdd vdd nmos L=40e-9 W=180e-9
m719 net07593 net07580 vdd vdd nmos L=40e-9 W=180e-9
m716 net07580 c28 vdd vdd nmos L=40e-9 W=180e-9
m715 net07580 net07576 vdd vdd nmos L=40e-9 W=180e-9
m712 net07513 net07507 vdd vdd nmos L=40e-9 W=180e-9
m711 net07513 net07494 vdd vdd nmos L=40e-9 W=180e-9
m710 net07546 net07527 vdd vdd nmos L=40e-9 W=180e-9
m709 net07546 net07540 vdd vdd nmos L=40e-9 W=180e-9
m708 net07358 net07340 vdd vdd nmos L=40e-9 W=180e-9
m707 net07358 net07352 vdd vdd nmos L=40e-9 W=180e-9
m706 net07389 net07370 vdd vdd nmos L=40e-9 W=180e-9
m705 net07389 net07383 vdd vdd nmos L=40e-9 W=180e-9
m704 net07420 net07414 vdd vdd nmos L=40e-9 W=180e-9
m703 net07420 net07401 vdd vdd nmos L=40e-9 W=180e-9
m702 net07451 net07432 vdd vdd nmos L=40e-9 W=180e-9
m701 net07451 net07445 vdd vdd nmos L=40e-9 W=180e-9
m700 net07482 net07476 vdd vdd nmos L=40e-9 W=180e-9
m699 net07482 net07463 vdd vdd nmos L=40e-9 W=180e-9
m698 net07507 c26 vdd vdd nmos L=40e-9 W=180e-9
m697 net07540 c27 vdd vdd nmos L=40e-9 W=180e-9
m696 net07572 c28 vdd vdd nmos L=40e-9 W=180e-9
m695 net07352 c22 vdd vdd nmos L=40e-9 W=180e-9
m694 net07383 c23 vdd vdd nmos L=40e-9 W=180e-9
m693 net07414 c24 vdd vdd nmos L=40e-9 W=180e-9
m692 net07445 net08819 vdd vdd nmos L=40e-9 W=180e-9
m691 net07476 c25 vdd vdd nmos L=40e-9 W=180e-9
m668 net07527 net07513 vdd vdd nmos L=40e-9 W=180e-9
m667 net07527 net07516 vdd vdd nmos L=40e-9 W=180e-9
m666 net07559 net07548 vdd vdd nmos L=40e-9 W=180e-9
m665 net07559 net07546 vdd vdd nmos L=40e-9 W=180e-9
m664 net07370 net07360 vdd vdd nmos L=40e-9 W=180e-9
m663 net07370 net07358 vdd vdd nmos L=40e-9 W=180e-9
m662 net07401 net07391 vdd vdd nmos L=40e-9 W=180e-9
m661 net07401 net07389 vdd vdd nmos L=40e-9 W=180e-9
m660 net07432 net07420 vdd vdd nmos L=40e-9 W=180e-9
m659 net07432 net07422 vdd vdd nmos L=40e-9 W=180e-9
m658 net07463 net07453 vdd vdd nmos L=40e-9 W=180e-9
m657 net07463 net07451 vdd vdd nmos L=40e-9 W=180e-9
m656 net07494 net07482 vdd vdd nmos L=40e-9 W=180e-9
m655 net07494 net07484 vdd vdd nmos L=40e-9 W=180e-9
m640 net07516 c26 vdd vdd nmos L=40e-9 W=180e-9
m639 net07516 net07511 vdd vdd nmos L=40e-9 W=180e-9
m638 net07548 net07544 vdd vdd nmos L=40e-9 W=180e-9
m637 net07548 c27 vdd vdd nmos L=40e-9 W=180e-9
m636 net07360 net07356 vdd vdd nmos L=40e-9 W=180e-9
m635 net07360 c22 vdd vdd nmos L=40e-9 W=180e-9
m634 net07391 net07387 vdd vdd nmos L=40e-9 W=180e-9
m633 net07391 c23 vdd vdd nmos L=40e-9 W=180e-9
m632 net07422 c24 vdd vdd nmos L=40e-9 W=180e-9
m631 net07422 net07418 vdd vdd nmos L=40e-9 W=180e-9
m630 net07453 net07449 vdd vdd nmos L=40e-9 W=180e-9
m629 net07453 net08819 vdd vdd nmos L=40e-9 W=180e-9
m628 net07484 c25 vdd vdd nmos L=40e-9 W=180e-9
m627 net07484 net07480 vdd vdd nmos L=40e-9 W=180e-9
m612 net07325 net07306 vdd vdd nmos L=40e-9 W=180e-9
m611 net07325 net07319 vdd vdd nmos L=40e-9 W=180e-9
m610 net07294 net07288 vdd vdd nmos L=40e-9 W=180e-9
m609 net07294 net07275 vdd vdd nmos L=40e-9 W=180e-9
m608 net07263 net07244 vdd vdd nmos L=40e-9 W=180e-9
m607 net07263 net07257 vdd vdd nmos L=40e-9 W=180e-9
m606 net07231 net07212 vdd vdd nmos L=40e-9 W=180e-9
m605 net07231 net07225 vdd vdd nmos L=40e-9 W=180e-9
m604 net07200 net07194 vdd vdd nmos L=40e-9 W=180e-9
m603 net07200 net07181 vdd vdd nmos L=40e-9 W=180e-9
m602 net07169 net07150 vdd vdd nmos L=40e-9 W=180e-9
m601 net07169 net07163 vdd vdd nmos L=40e-9 W=180e-9
m600 net07138 net07132 vdd vdd nmos L=40e-9 W=180e-9
m599 net07138 net07119 vdd vdd nmos L=40e-9 W=180e-9
m598 net07107 net07101 vdd vdd nmos L=40e-9 W=180e-9
m597 net07107 net07089 vdd vdd nmos L=40e-9 W=180e-9
m596 net07319 c21 vdd vdd nmos L=40e-9 W=180e-9
m595 net07288 c20 vdd vdd nmos L=40e-9 W=180e-9
m594 net07257 c19 vdd vdd nmos L=40e-9 W=180e-9
m593 net07225 c18 vdd vdd nmos L=40e-9 W=180e-9
m592 net07194 c17 vdd vdd nmos L=40e-9 W=180e-9
m591 net07163 net08803 vdd vdd nmos L=40e-9 W=180e-9
m590 net07132 c16 vdd vdd nmos L=40e-9 W=180e-9
m589 net07101 c15 vdd vdd nmos L=40e-9 W=180e-9
m569 net07340 net07327 vdd vdd nmos L=40e-9 W=180e-9
m568 net07340 net07325 vdd vdd nmos L=40e-9 W=180e-9
m567 net07306 net07294 vdd vdd nmos L=40e-9 W=180e-9
m566 net07306 net07296 vdd vdd nmos L=40e-9 W=180e-9
m565 net07275 net07265 vdd vdd nmos L=40e-9 W=180e-9
m564 net07275 net07263 vdd vdd nmos L=40e-9 W=180e-9
m558 net07244 net07234 vdd vdd nmos L=40e-9 W=180e-9
m557 net07244 net07231 vdd vdd nmos L=40e-9 W=180e-9
m556 net07212 net07200 vdd vdd nmos L=40e-9 W=180e-9
m555 net07212 net07202 vdd vdd nmos L=40e-9 W=180e-9
m554 net07181 net07171 vdd vdd nmos L=40e-9 W=180e-9
m553 net07181 net07169 vdd vdd nmos L=40e-9 W=180e-9
m552 net07150 net07138 vdd vdd nmos L=40e-9 W=180e-9
m551 net07150 net07140 vdd vdd nmos L=40e-9 W=180e-9
m550 net07119 net07107 vdd vdd nmos L=40e-9 W=180e-9
m549 net07119 net07109 vdd vdd nmos L=40e-9 W=180e-9
m532 net07327 net07323 vdd vdd nmos L=40e-9 W=180e-9
m531 net07327 c21 vdd vdd nmos L=40e-9 W=180e-9
m530 net07296 c20 vdd vdd nmos L=40e-9 W=180e-9
m529 net07296 net07292 vdd vdd nmos L=40e-9 W=180e-9
m528 net07265 net07261 vdd vdd nmos L=40e-9 W=180e-9
m527 net07265 c19 vdd vdd nmos L=40e-9 W=180e-9
m526 net07234 net07229 vdd vdd nmos L=40e-9 W=180e-9
m525 net07234 c18 vdd vdd nmos L=40e-9 W=180e-9
m524 net07202 c17 vdd vdd nmos L=40e-9 W=180e-9
m523 net07202 net07198 vdd vdd nmos L=40e-9 W=180e-9
m522 net07171 net07167 vdd vdd nmos L=40e-9 W=180e-9
m521 net07171 net08803 vdd vdd nmos L=40e-9 W=180e-9
m520 net07140 c16 vdd vdd nmos L=40e-9 W=180e-9
m519 net07140 net07136 vdd vdd nmos L=40e-9 W=180e-9
m518 net07109 c15 vdd vdd nmos L=40e-9 W=180e-9
m517 net07109 net07105 vdd vdd nmos L=40e-9 W=180e-9
m500 net07076 net07067 vdd vdd nmos L=40e-9 W=180e-9
m499 net07041 net07033 vdd vdd nmos L=40e-9 W=180e-9
m498 net07041 net07034 vdd vdd nmos L=40e-9 W=180e-9
m497 net07076 net07068 vdd vdd nmos L=40e-9 W=180e-9
m496 net07007 net06998 vdd vdd nmos L=40e-9 W=180e-9
m495 net07007 net06997 vdd vdd nmos L=40e-9 W=180e-9
m494 net07067 c14 vdd vdd nmos L=40e-9 W=180e-9
m493 net07033 c13 vdd vdd nmos L=40e-9 W=180e-9
m484 net07105 net07076 vdd vdd nmos L=40e-9 W=180e-9
m483 net07068 net07041 vdd vdd nmos L=40e-9 W=180e-9
m482 net07068 net07044 vdd vdd nmos L=40e-9 W=180e-9
m481 net07034 net07010 vdd vdd nmos L=40e-9 W=180e-9
m480 net07034 net07007 vdd vdd nmos L=40e-9 W=180e-9
m479 net07105 net07079 vdd vdd nmos L=40e-9 W=180e-9
m478 net06973 net06966 vdd vdd nmos L=40e-9 W=180e-9
m477 net06942 net06935 vdd vdd nmos L=40e-9 W=180e-9
m476 net06942 net06936 vdd vdd nmos L=40e-9 W=180e-9
m475 net06973 net06967 vdd vdd nmos L=40e-9 W=180e-9
m474 net06997 c12 vdd vdd nmos L=40e-9 W=180e-9
m473 net06966 c11 vdd vdd nmos L=40e-9 W=180e-9
m472 net06935 c10 vdd vdd nmos L=40e-9 W=180e-9
m464 net06998 net06975 vdd vdd nmos L=40e-9 W=180e-9
m463 net06998 net06973 vdd vdd nmos L=40e-9 W=180e-9
m462 net06967 net06942 vdd vdd nmos L=40e-9 W=180e-9
m461 net06967 net06944 vdd vdd nmos L=40e-9 W=180e-9
m460 net06936 net06913 vdd vdd nmos L=40e-9 W=180e-9
m459 net06936 net06911 vdd vdd nmos L=40e-9 W=180e-9
m458 net06911 net06905 vdd vdd nmos L=40e-9 W=180e-9
m457 net06911 net06904 vdd vdd nmos L=40e-9 W=180e-9
m456 net06880 net06873 vdd vdd nmos L=40e-9 W=180e-9
m455 net06880 net06874 vdd vdd nmos L=40e-9 W=180e-9
m454 net06849 net06842 vdd vdd nmos L=40e-9 W=180e-9
m453 net06849 net0988 vdd vdd nmos L=40e-9 W=180e-9
m452 net06904 c9 vdd vdd nmos L=40e-9 W=180e-9
m451 net06873 net08787 vdd vdd nmos L=40e-9 W=180e-9
m450 net06842 c8 vdd vdd nmos L=40e-9 W=180e-9
m440 net06905 net06880 vdd vdd nmos L=40e-9 W=180e-9
m439 net06905 net06882 vdd vdd nmos L=40e-9 W=180e-9
m438 net06874 net06849 vdd vdd nmos L=40e-9 W=180e-9
m437 net06874 net06851 vdd vdd nmos L=40e-9 W=180e-9
m430 net07079 net07051 vdd vdd nmos L=40e-9 W=180e-9
m429 net07079 c14 vdd vdd nmos L=40e-9 W=180e-9
m428 net07044 c13 vdd vdd nmos L=40e-9 W=180e-9
m427 net07044 net07017 vdd vdd nmos L=40e-9 W=180e-9
m426 net07010 net06981 vdd vdd nmos L=40e-9 W=180e-9
m425 net07010 c12 vdd vdd nmos L=40e-9 W=180e-9
m412 net06975 net06950 vdd vdd nmos L=40e-9 W=180e-9
m411 net06975 c11 vdd vdd nmos L=40e-9 W=180e-9
m410 net06944 c10 vdd vdd nmos L=40e-9 W=180e-9
m409 net06944 net06919 vdd vdd nmos L=40e-9 W=180e-9
m400 net06913 net06888 vdd vdd nmos L=40e-9 W=180e-9
m399 net06913 c9 vdd vdd nmos L=40e-9 W=180e-9
m398 net06882 net08787 vdd vdd nmos L=40e-9 W=180e-9
m397 net06882 net06857 vdd vdd nmos L=40e-9 W=180e-9
m396 net06851 c8 vdd vdd nmos L=40e-9 W=180e-9
m395 net06851 net0955 vdd vdd nmos L=40e-9 W=180e-9
m388 net07071 net07051 vdd vdd nmos L=40e-9 W=180e-9
m387 net07071 net07064 vdd vdd nmos L=40e-9 W=180e-9
m386 net07036 net07030 vdd vdd nmos L=40e-9 W=180e-9
m385 net07036 net07017 vdd vdd nmos L=40e-9 W=180e-9
m384 net07001 net06981 vdd vdd nmos L=40e-9 W=180e-9
m383 net07001 net06994 vdd vdd nmos L=40e-9 W=180e-9
m382 net07064 c14 vdd vdd nmos L=40e-9 W=180e-9
m381 net07030 c13 vdd vdd nmos L=40e-9 W=180e-9
m372 net07089 net07074 vdd vdd nmos L=40e-9 W=180e-9
m371 net07089 net07071 vdd vdd nmos L=40e-9 W=180e-9
m370 net07051 net07036 vdd vdd nmos L=40e-9 W=180e-9
m369 net07051 net07039 vdd vdd nmos L=40e-9 W=180e-9
m368 net07017 net07004 vdd vdd nmos L=40e-9 W=180e-9
m367 net07017 net07001 vdd vdd nmos L=40e-9 W=180e-9
m360 net07074 net07068 vdd vdd nmos L=40e-9 W=180e-9
m359 net07074 c14 vdd vdd nmos L=40e-9 W=180e-9
m358 net07039 c13 vdd vdd nmos L=40e-9 W=180e-9
m357 net07039 net07034 vdd vdd nmos L=40e-9 W=180e-9
m356 net07004 net06998 vdd vdd nmos L=40e-9 W=180e-9
m355 net07004 c12 vdd vdd nmos L=40e-9 W=180e-9
m348 net06969 net06950 vdd vdd nmos L=40e-9 W=180e-9
m347 net06969 net06963 vdd vdd nmos L=40e-9 W=180e-9
m346 net06938 net06932 vdd vdd nmos L=40e-9 W=180e-9
m345 net06938 net06919 vdd vdd nmos L=40e-9 W=180e-9
m344 net06994 c12 vdd vdd nmos L=40e-9 W=180e-9
m343 net06963 c11 vdd vdd nmos L=40e-9 W=180e-9
m342 net06932 c10 vdd vdd nmos L=40e-9 W=180e-9
m334 net06981 net06971 vdd vdd nmos L=40e-9 W=180e-9
m333 net06981 net06969 vdd vdd nmos L=40e-9 W=180e-9
m332 net06950 net06938 vdd vdd nmos L=40e-9 W=180e-9
m331 net06950 net06940 vdd vdd nmos L=40e-9 W=180e-9
m330 net06919 net06909 vdd vdd nmos L=40e-9 W=180e-9
m329 net06919 net06907 vdd vdd nmos L=40e-9 W=180e-9
m322 net06971 net06967 vdd vdd nmos L=40e-9 W=180e-9
m321 net06971 c11 vdd vdd nmos L=40e-9 W=180e-9
m320 net06940 c10 vdd vdd nmos L=40e-9 W=180e-9
m319 net06940 net06936 vdd vdd nmos L=40e-9 W=180e-9
m314 net06907 net06888 vdd vdd nmos L=40e-9 W=180e-9
m313 net06907 net06901 vdd vdd nmos L=40e-9 W=180e-9
m312 net06876 net06870 vdd vdd nmos L=40e-9 W=180e-9
m311 net06876 net06857 vdd vdd nmos L=40e-9 W=180e-9
m310 net06845 net06839 vdd vdd nmos L=40e-9 W=180e-9
m309 net06845 net0955 vdd vdd nmos L=40e-9 W=180e-9
m308 net06901 c9 vdd vdd nmos L=40e-9 W=180e-9
m307 net06870 net08787 vdd vdd nmos L=40e-9 W=180e-9
m306 net06839 c8 vdd vdd nmos L=40e-9 W=180e-9
m296 net06888 net06876 vdd vdd nmos L=40e-9 W=180e-9
m295 net06888 net06878 vdd vdd nmos L=40e-9 W=180e-9
m294 net06857 net06845 vdd vdd nmos L=40e-9 W=180e-9
m293 net06857 net06847 vdd vdd nmos L=40e-9 W=180e-9
m288 net06909 net06905 vdd vdd nmos L=40e-9 W=180e-9
m287 net06909 c9 vdd vdd nmos L=40e-9 W=180e-9
m286 net06878 net08787 vdd vdd nmos L=40e-9 W=180e-9
m285 net06878 net06874 vdd vdd nmos L=40e-9 W=180e-9
m284 net06847 c8 vdd vdd nmos L=40e-9 W=180e-9
m283 net06847 net0988 vdd vdd nmos L=40e-9 W=180e-9
m250 net0947 net0940 vdd vdd nmos L=40e-9 W=180e-9
m249 net0947 net0941 vdd vdd nmos L=40e-9 W=180e-9
m247 net0916 net0910 vdd vdd nmos L=40e-9 W=180e-9
m246 net0916 net0909 vdd vdd nmos L=40e-9 W=180e-9
m244 net0940 c7 vdd vdd nmos L=40e-9 W=180e-9
m243 net0909 c6 vdd vdd nmos L=40e-9 W=180e-9
m232 net0988 net0947 vdd vdd nmos L=40e-9 W=180e-9
m231 net0988 net0949 vdd vdd nmos L=40e-9 W=180e-9
m230 net0941 net0918 vdd vdd nmos L=40e-9 W=180e-9
m229 net0941 net0916 vdd vdd nmos L=40e-9 W=180e-9
m220 net0949 c7 vdd vdd nmos L=40e-9 W=180e-9
m219 net0949 net0924 vdd vdd nmos L=40e-9 W=180e-9
m218 net0918 net0893 vdd vdd nmos L=40e-9 W=180e-9
m217 net0918 c6 vdd vdd nmos L=40e-9 W=180e-9
m208 net0943 net0937 vdd vdd nmos L=40e-9 W=180e-9
m207 net0943 net0924 vdd vdd nmos L=40e-9 W=180e-9
m206 net0912 net0893 vdd vdd nmos L=40e-9 W=180e-9
m205 net0912 net0906 vdd vdd nmos L=40e-9 W=180e-9
m203 net0937 c7 vdd vdd nmos L=40e-9 W=180e-9
m202 net0906 c6 vdd vdd nmos L=40e-9 W=180e-9
m190 net0955 net0943 vdd vdd nmos L=40e-9 W=180e-9
m189 net0955 net0945 vdd vdd nmos L=40e-9 W=180e-9
m188 net0924 net0914 vdd vdd nmos L=40e-9 W=180e-9
m187 net0924 net0912 vdd vdd nmos L=40e-9 W=180e-9
m178 net0945 c7 vdd vdd nmos L=40e-9 W=180e-9
m177 net0945 net0941 vdd vdd nmos L=40e-9 W=180e-9
m176 net0914 net0910 vdd vdd nmos L=40e-9 W=180e-9
m175 net0914 c6 vdd vdd nmos L=40e-9 W=180e-9
m167 net0885 net0879 vdd vdd nmos L=40e-9 W=180e-9
m166 net0885 net0878 vdd vdd nmos L=40e-9 W=180e-9
m165 net0854 net0847 vdd vdd nmos L=40e-9 W=180e-9
m164 net0854 net0848 vdd vdd nmos L=40e-9 W=180e-9
m163 net0878 c5 vdd vdd nmos L=40e-9 W=180e-9
m162 net0847 c4 vdd vdd nmos L=40e-9 W=180e-9
m155 net0910 net0885 vdd vdd nmos L=40e-9 W=180e-9
m154 net0879 net0854 vdd vdd nmos L=40e-9 W=180e-9
m153 net0879 net0856 vdd vdd nmos L=40e-9 W=180e-9
m148 net0887 net0862 vdd vdd nmos L=40e-9 W=180e-9
m147 net0887 c5 vdd vdd nmos L=40e-9 W=180e-9
m146 net0856 c4 vdd vdd nmos L=40e-9 W=180e-9
m145 net0856 net0831 vdd vdd nmos L=40e-9 W=180e-9
m140 net0881 net0862 vdd vdd nmos L=40e-9 W=180e-9
m139 net0881 net0875 vdd vdd nmos L=40e-9 W=180e-9
m138 net0850 net0844 vdd vdd nmos L=40e-9 W=180e-9
m137 net0850 net0831 vdd vdd nmos L=40e-9 W=180e-9
m136 net0875 c5 vdd vdd nmos L=40e-9 W=180e-9
m135 net0844 c4 vdd vdd nmos L=40e-9 W=180e-9
m128 net0893 net0883 vdd vdd nmos L=40e-9 W=180e-9
m127 net0893 net0881 vdd vdd nmos L=40e-9 W=180e-9
m126 net0862 net0850 vdd vdd nmos L=40e-9 W=180e-9
m125 net0862 net0852 vdd vdd nmos L=40e-9 W=180e-9
m120 net0883 net0879 vdd vdd nmos L=40e-9 W=180e-9
m119 net0883 c5 vdd vdd nmos L=40e-9 W=180e-9
m118 net0852 c4 vdd vdd nmos L=40e-9 W=180e-9
m117 net0852 net0848 vdd vdd nmos L=40e-9 W=180e-9
m112 net0910 net0887 vdd vdd nmos L=40e-9 W=180e-9
m111 net0823 net0816 vdd vdd nmos L=40e-9 W=180e-9
m110 net0823 net0200 vdd vdd nmos L=40e-9 W=180e-9
m109 net0816 c3 vdd vdd nmos L=40e-9 W=180e-9
m105 net0848 net0823 vdd vdd nmos L=40e-9 W=180e-9
m104 net0848 net0825 vdd vdd nmos L=40e-9 W=180e-9
m101 net0825 c3 vdd vdd nmos L=40e-9 W=180e-9
m100 net0825 net0198 vdd vdd nmos L=40e-9 W=180e-9
m97 net0819 net0813 vdd vdd nmos L=40e-9 W=180e-9
m96 net0819 net0198 vdd vdd nmos L=40e-9 W=180e-9
m95 net0813 c3 vdd vdd nmos L=40e-9 W=180e-9
m91 net0831 net0819 vdd vdd nmos L=40e-9 W=180e-9
m90 net0831 net0821 vdd vdd nmos L=40e-9 W=180e-9
m87 net0821 c3 vdd vdd nmos L=40e-9 W=180e-9
m86 net0821 net0200 vdd vdd nmos L=40e-9 W=180e-9
m83 net0190 net0183 vdd vdd nmos L=40e-9 W=180e-9
m82 net0190 net55 vdd vdd nmos L=40e-9 W=180e-9
m81 net0183 c2 vdd vdd nmos L=40e-9 W=180e-9
m77 net0200 net0190 vdd vdd nmos L=40e-9 W=180e-9
m76 net0200 net0192 vdd vdd nmos L=40e-9 W=180e-9
m73 net0192 c2 vdd vdd nmos L=40e-9 W=180e-9
m72 net0192 net51 vdd vdd nmos L=40e-9 W=180e-9
m69 net0186 net0180 vdd vdd nmos L=40e-9 W=180e-9
m68 net0186 net51 vdd vdd nmos L=40e-9 W=180e-9
m67 net0180 c2 vdd vdd nmos L=40e-9 W=180e-9
m63 net0198 net0186 vdd vdd nmos L=40e-9 W=180e-9
m62 net0198 net0188 vdd vdd nmos L=40e-9 W=180e-9
m59 net0188 c2 vdd vdd nmos L=40e-9 W=180e-9
m58 net0188 net55 vdd vdd nmos L=40e-9 W=180e-9
m25 net51 net28 vdd vdd nmos L=40e-9 W=180e-9
m24 net51 net32 vdd vdd nmos L=40e-9 W=180e-9
m21 net32 c1 vdd vdd nmos L=40e-9 W=180e-9
m20 net32 start1 vdd vdd nmos L=40e-9 W=180e-9
m18 net19 c1 vdd vdd nmos L=40e-9 W=180e-9
m15 net28 net19 vdd vdd nmos L=40e-9 W=180e-9
m14 net28 start2 vdd vdd nmos L=40e-9 W=180e-9
m11 net55 net36 vdd vdd nmos L=40e-9 W=180e-9
m10 net55 net39 vdd vdd nmos L=40e-9 W=180e-9
m7 net39 c1 vdd vdd nmos L=40e-9 W=180e-9
m6 net39 start2 vdd vdd nmos L=40e-9 W=180e-9
m4 net22 c1 vdd vdd nmos L=40e-9 W=180e-9
m3 net36 start1 vdd vdd nmos L=40e-9 W=180e-9
m1 net36 net22 vdd vdd nmos L=40e-9 W=180e-9
m2072 net04309 net04302 net06154 vss nmos L=40e-9 W=90e-9
m2071 net04489 net04482 net06148 vss nmos L=40e-9 W=90e-9
m2070 net04519 net04512 net06147 vss nmos L=40e-9 W=90e-9
m2069 net04459 net04452 net06149 vss nmos L=40e-9 W=90e-9
m2068 net04429 net04422 net06150 vss nmos L=40e-9 W=90e-9
m2067 net04399 net04392 net06151 vss nmos L=40e-9 W=90e-9
m2066 net04369 net04362 net06152 vss nmos L=40e-9 W=90e-9
m2065 net04339 net04332 net06153 vss nmos L=40e-9 W=90e-9
m2064 net04302 c57 vss vss nmos L=40e-9 W=90e-9
m2063 net04482 c63 vss vss nmos L=40e-9 W=90e-9
m2062 net04512 c64 vss vss nmos L=40e-9 W=90e-9
m2061 net04452 c62 vss vss nmos L=40e-9 W=90e-9
m2060 net04422 c61 vss vss nmos L=40e-9 W=90e-9
m2059 net04392 c60 vss vss nmos L=40e-9 W=90e-9
m2058 net04362 c59 vss vss nmos L=40e-9 W=90e-9
m2057 net04332 c58 vss vss nmos L=40e-9 W=90e-9
m2056 net06154 net03543 vss vss nmos L=40e-9 W=90e-9
m2053 net06148 net04483 vss vss nmos L=40e-9 W=90e-9
m2052 net06147 net04513 vss vss nmos L=40e-9 W=90e-9
m2049 net06149 net04453 vss vss nmos L=40e-9 W=90e-9
m2048 net06150 net04423 vss vss nmos L=40e-9 W=90e-9
m2047 net06151 net04393 vss vss nmos L=40e-9 W=90e-9
m2044 net06152 net04363 vss vss nmos L=40e-9 W=90e-9
m2043 net06153 net04333 vss vss nmos L=40e-9 W=90e-9
m2032 net04333 net04309 net06162 vss nmos L=40e-9 W=90e-9
m2031 net04513 net04489 net06156 vss nmos L=40e-9 W=90e-9
m2030 net04550 net04519 net06155 vss nmos L=40e-9 W=90e-9
m2029 net04483 net04459 net06157 vss nmos L=40e-9 W=90e-9
m2028 net04453 net04429 net06158 vss nmos L=40e-9 W=90e-9
m2027 net04423 net04399 net06159 vss nmos L=40e-9 W=90e-9
m2026 net04393 net04369 net06160 vss nmos L=40e-9 W=90e-9
m2025 net04363 net04339 net06161 vss nmos L=40e-9 W=90e-9
m2024 net06162 net04311 vss vss nmos L=40e-9 W=90e-9
m2023 net06156 net04491 vss vss nmos L=40e-9 W=90e-9
m2022 net06155 net04521 vss vss nmos L=40e-9 W=90e-9
m2019 net06157 net04461 vss vss nmos L=40e-9 W=90e-9
m2018 net06158 net04431 vss vss nmos L=40e-9 W=90e-9
m2017 net06159 net04401 vss vss nmos L=40e-9 W=90e-9
m2016 net06160 net04371 vss vss nmos L=40e-9 W=90e-9
m2015 net06161 net04341 vss vss nmos L=40e-9 W=90e-9
m2000 net04311 c57 net06170 vss nmos L=40e-9 W=90e-9
m1999 net04491 c63 net06164 vss nmos L=40e-9 W=90e-9
m1998 net04521 c64 net06163 vss nmos L=40e-9 W=90e-9
m1997 net04461 c62 net06165 vss nmos L=40e-9 W=90e-9
m1996 net04431 c61 net06166 vss nmos L=40e-9 W=90e-9
m1995 net04401 c60 net06167 vss nmos L=40e-9 W=90e-9
m1994 net04371 c59 net06168 vss nmos L=40e-9 W=90e-9
m1993 net04341 c58 net06169 vss nmos L=40e-9 W=90e-9
m1992 net06170 net08593 vss vss nmos L=40e-9 W=90e-9
m1991 net06164 net04467 vss vss nmos L=40e-9 W=90e-9
m1990 net06163 net04497 vss vss nmos L=40e-9 W=90e-9
m1989 net06165 net04437 vss vss nmos L=40e-9 W=90e-9
m1988 net06166 net04407 vss vss nmos L=40e-9 W=90e-9
m1987 net06167 net04377 vss vss nmos L=40e-9 W=90e-9
m1986 net06168 net04347 vss vss nmos L=40e-9 W=90e-9
m1985 net06169 net04317 vss vss nmos L=40e-9 W=90e-9
m1960 net04305 net04299 net06171 vss nmos L=40e-9 W=90e-9
m1959 net04485 net04479 net06173 vss nmos L=40e-9 W=90e-9
m1958 net04515 net04509 net06172 vss nmos L=40e-9 W=90e-9
m1957 net04395 net04389 net06176 vss nmos L=40e-9 W=90e-9
m1956 net04425 net04419 net06175 vss nmos L=40e-9 W=90e-9
m1955 net04455 net04449 net06174 vss nmos L=40e-9 W=90e-9
m1954 net04335 net04329 net06178 vss nmos L=40e-9 W=90e-9
m1953 net04365 net04359 net06177 vss nmos L=40e-9 W=90e-9
m1952 net04299 c57 vss vss nmos L=40e-9 W=90e-9
m1951 net04479 c63 vss vss nmos L=40e-9 W=90e-9
m1950 net04509 c64 vss vss nmos L=40e-9 W=90e-9
m1949 net04389 c60 vss vss nmos L=40e-9 W=90e-9
m1948 net04419 c61 vss vss nmos L=40e-9 W=90e-9
m1947 net04449 c62 vss vss nmos L=40e-9 W=90e-9
m1946 net04329 c58 vss vss nmos L=40e-9 W=90e-9
m1945 net04359 c59 vss vss nmos L=40e-9 W=90e-9
m1944 net06171 net08593 vss vss nmos L=40e-9 W=90e-9
m1941 net06173 net04467 vss vss nmos L=40e-9 W=90e-9
m1940 net06172 net04497 vss vss nmos L=40e-9 W=90e-9
m1939 net06176 net04377 vss vss nmos L=40e-9 W=90e-9
m1938 net06175 net04407 vss vss nmos L=40e-9 W=90e-9
m1937 net06174 net04437 vss vss nmos L=40e-9 W=90e-9
m1932 net06178 net04317 vss vss nmos L=40e-9 W=90e-9
m1931 net06177 net04347 vss vss nmos L=40e-9 W=90e-9
m1920 net04317 net04305 net06179 vss nmos L=40e-9 W=90e-9
m1919 net04497 net04485 net06181 vss nmos L=40e-9 W=90e-9
m1918 net04530 net04515 net06180 vss nmos L=40e-9 W=90e-9
m1917 net04407 net04395 net06184 vss nmos L=40e-9 W=90e-9
m1916 net04437 net04425 net06183 vss nmos L=40e-9 W=90e-9
m1915 net04467 net04455 net06182 vss nmos L=40e-9 W=90e-9
m1914 net04347 net04335 net06186 vss nmos L=40e-9 W=90e-9
m1913 net04377 net04365 net06185 vss nmos L=40e-9 W=90e-9
m1912 net06179 net04307 vss vss nmos L=40e-9 W=90e-9
m1911 net06181 net04487 vss vss nmos L=40e-9 W=90e-9
m1910 net06180 net04517 vss vss nmos L=40e-9 W=90e-9
m1907 net06184 net04397 vss vss nmos L=40e-9 W=90e-9
m1906 net06183 net04427 vss vss nmos L=40e-9 W=90e-9
m1905 net06182 net04457 vss vss nmos L=40e-9 W=90e-9
m1904 net06186 net04337 vss vss nmos L=40e-9 W=90e-9
m1903 net06185 net04367 vss vss nmos L=40e-9 W=90e-9
m1888 net04307 c57 net06194 vss nmos L=40e-9 W=90e-9
m1887 net04487 c63 net06188 vss nmos L=40e-9 W=90e-9
m1886 net04517 c64 net06187 vss nmos L=40e-9 W=90e-9
m1885 net04397 c60 net06191 vss nmos L=40e-9 W=90e-9
m1884 net04427 c61 net06190 vss nmos L=40e-9 W=90e-9
m1883 net04457 c62 net06189 vss nmos L=40e-9 W=90e-9
m1882 net04337 c58 net06193 vss nmos L=40e-9 W=90e-9
m1881 net04367 c59 net06192 vss nmos L=40e-9 W=90e-9
m1880 net06194 net03543 vss vss nmos L=40e-9 W=90e-9
m1879 net06188 net04483 vss vss nmos L=40e-9 W=90e-9
m1878 net06187 net04513 vss vss nmos L=40e-9 W=90e-9
m1877 net06191 net04393 vss vss nmos L=40e-9 W=90e-9
m1876 net06190 net04423 vss vss nmos L=40e-9 W=90e-9
m1875 net06189 net04453 vss vss nmos L=40e-9 W=90e-9
m1874 net06192 net04363 vss vss nmos L=40e-9 W=90e-9
m1873 net06193 net04333 vss vss nmos L=40e-9 W=90e-9
m1869 net03549 net03542 net05100 vss nmos L=40e-9 W=90e-9
m1868 net03542 net05098 vss vss nmos L=40e-9 W=90e-9
m1867 net05100 net04550 vss vss nmos L=40e-9 W=90e-9
m1864 net03559 net03549 net05101 vss nmos L=40e-9 W=90e-9
m1863 net05101 net03551 vss vss nmos L=40e-9 W=90e-9
m1860 net03551 net05098 net05102 vss nmos L=40e-9 W=90e-9
m1859 net05102 net04530 vss vss nmos L=40e-9 W=90e-9
m1855 net03545 net03539 net05103 vss nmos L=40e-9 W=90e-9
m1854 net03539 net05098 vss vss nmos L=40e-9 W=90e-9
m1853 net05103 net04530 vss vss nmos L=40e-9 W=90e-9
m1850 net03557 net03545 net05104 vss nmos L=40e-9 W=90e-9
m1849 net05104 net03547 vss vss nmos L=40e-9 W=90e-9
m1846 net03547 net05098 net05105 vss nmos L=40e-9 W=90e-9
m1845 net05105 net04550 vss vss nmos L=40e-9 W=90e-9
m1838 net08551 net08544 net08902 vss nmos L=40e-9 W=90e-9
m1837 net08582 net08575 net08901 vss nmos L=40e-9 W=90e-9
m1836 net08544 c56 vss vss nmos L=40e-9 W=90e-9
m1835 net08575 net08884 vss vss nmos L=40e-9 W=90e-9
m1834 net08902 net08545 vss vss nmos L=40e-9 W=90e-9
m1833 net08901 net08576 vss vss nmos L=40e-9 W=90e-9
m1828 net08576 net08551 net08934 vss nmos L=40e-9 W=90e-9
m1827 net03543 net08582 net08933 vss nmos L=40e-9 W=90e-9
m1781 net08270 net08263 net08911 vss nmos L=40e-9 W=90e-9
m1780 net08301 net08294 net08910 vss nmos L=40e-9 W=90e-9
m1779 net08332 net08325 net08909 vss nmos L=40e-9 W=90e-9
m1778 net08115 net08108 net08916 vss nmos L=40e-9 W=90e-9
m1777 net08146 net08139 net08915 vss nmos L=40e-9 W=90e-9
m1776 net08177 net08170 net08914 vss nmos L=40e-9 W=90e-9
m1775 net08208 net08201 net08913 vss nmos L=40e-9 W=90e-9
m1774 net08239 net08232 net08912 vss nmos L=40e-9 W=90e-9
m1773 net08082 net08075 net08917 vss nmos L=40e-9 W=90e-9
m1772 net08520 net08513 net08903 vss nmos L=40e-9 W=90e-9
m1771 net08365 net08358 net08908 vss nmos L=40e-9 W=90e-9
m1770 net08396 net08389 net08907 vss nmos L=40e-9 W=90e-9
m1769 net08427 net08420 net08906 vss nmos L=40e-9 W=90e-9
m1768 net08458 net08451 net08905 vss nmos L=40e-9 W=90e-9
m1767 net08489 net08482 net08904 vss nmos L=40e-9 W=90e-9
m1766 net08263 c48 vss vss nmos L=40e-9 W=90e-9
m1765 net08294 net08868 vss vss nmos L=40e-9 W=90e-9
m1764 net08325 c49 vss vss nmos L=40e-9 W=90e-9
m1763 net08108 c43 vss vss nmos L=40e-9 W=90e-9
m1762 net08139 c44 vss vss nmos L=40e-9 W=90e-9
m1761 net08170 c45 vss vss nmos L=40e-9 W=90e-9
m1760 net08201 c46 vss vss nmos L=40e-9 W=90e-9
m1759 net08232 c47 vss vss nmos L=40e-9 W=90e-9
m1758 net08075 c42 vss vss nmos L=40e-9 W=90e-9
m1757 net08513 c55 vss vss nmos L=40e-9 W=90e-9
m1756 net08358 c50 vss vss nmos L=40e-9 W=90e-9
m1755 net08389 c51 vss vss nmos L=40e-9 W=90e-9
m1754 net08420 c52 vss vss nmos L=40e-9 W=90e-9
m1753 net08451 c53 vss vss nmos L=40e-9 W=90e-9
m1752 net08482 c54 vss vss nmos L=40e-9 W=90e-9
m1751 net08911 net08264 vss vss nmos L=40e-9 W=90e-9
m1750 net08910 net08295 vss vss nmos L=40e-9 W=90e-9
m1749 net08909 net08326 vss vss nmos L=40e-9 W=90e-9
m1748 net08916 net08109 vss vss nmos L=40e-9 W=90e-9
m1747 net08915 net08140 vss vss nmos L=40e-9 W=90e-9
m1746 net08914 net08171 vss vss nmos L=40e-9 W=90e-9
m1745 net08913 net08202 vss vss nmos L=40e-9 W=90e-9
m1744 net08912 net08233 vss vss nmos L=40e-9 W=90e-9
m1737 net08917 net08076 vss vss nmos L=40e-9 W=90e-9
m1724 net08903 net08514 vss vss nmos L=40e-9 W=90e-9
m1723 net08908 net08359 vss vss nmos L=40e-9 W=90e-9
m1722 net08907 net08390 vss vss nmos L=40e-9 W=90e-9
m1721 net08906 net08421 vss vss nmos L=40e-9 W=90e-9
m1720 net08905 net08452 vss vss nmos L=40e-9 W=90e-9
m1719 net08904 net08483 vss vss nmos L=40e-9 W=90e-9
m1706 net08295 net08270 net08943 vss nmos L=40e-9 W=90e-9
m1705 net08326 net08301 net08942 vss nmos L=40e-9 W=90e-9
m1704 net08359 net08332 net08941 vss nmos L=40e-9 W=90e-9
m1703 net08140 net08115 net08948 vss nmos L=40e-9 W=90e-9
m1702 net08171 net08146 net08947 vss nmos L=40e-9 W=90e-9
m1701 net08202 net08177 net08946 vss nmos L=40e-9 W=90e-9
m1700 net08233 net08208 net08945 vss nmos L=40e-9 W=90e-9
m1699 net08264 net08239 net08944 vss nmos L=40e-9 W=90e-9
m1698 net08109 net08082 net08949 vss nmos L=40e-9 W=90e-9
m1697 net08545 net08520 net08935 vss nmos L=40e-9 W=90e-9
m1696 net08390 net08365 net08940 vss nmos L=40e-9 W=90e-9
m1695 net08421 net08396 net08939 vss nmos L=40e-9 W=90e-9
m1694 net08452 net08427 net08938 vss nmos L=40e-9 W=90e-9
m1693 net08483 net08458 net08937 vss nmos L=40e-9 W=90e-9
m1692 net08514 net08489 net08936 vss nmos L=40e-9 W=90e-9
m1691 net08943 net08272 vss vss nmos L=40e-9 W=90e-9
m1690 net08942 net08303 vss vss nmos L=40e-9 W=90e-9
m1689 net08941 net08334 vss vss nmos L=40e-9 W=90e-9
m1643 net07832 net07825 net08925 vss nmos L=40e-9 W=90e-9
m1642 net07801 net07794 net08926 vss nmos L=40e-9 W=90e-9
m1641 net07770 net07763 net08927 vss nmos L=40e-9 W=90e-9
m1640 net07739 net07732 net08928 vss nmos L=40e-9 W=90e-9
m1639 net07708 net07701 net08929 vss nmos L=40e-9 W=90e-9
m1638 net07677 net07670 net08930 vss nmos L=40e-9 W=90e-9
m1637 net07646 net07639 net08931 vss nmos L=40e-9 W=90e-9
m1636 net07615 net07608 net08932 vss nmos L=40e-9 W=90e-9
m1635 net08051 net08044 net08918 vss nmos L=40e-9 W=90e-9
m1634 net08020 net08013 net08919 vss nmos L=40e-9 W=90e-9
m1633 net07989 net07982 net08920 vss nmos L=40e-9 W=90e-9
m1632 net07958 net07951 net08921 vss nmos L=40e-9 W=90e-9
m1631 net07927 net07920 net08922 vss nmos L=40e-9 W=90e-9
m1630 net07896 net07889 net08923 vss nmos L=40e-9 W=90e-9
m1629 net07865 net07858 net08924 vss nmos L=40e-9 W=90e-9
m1628 net07825 c35 vss vss nmos L=40e-9 W=90e-9
m1627 net07794 c34 vss vss nmos L=40e-9 W=90e-9
m1626 net07763 c33 vss vss nmos L=40e-9 W=90e-9
m1625 net07732 net08836 vss vss nmos L=40e-9 W=90e-9
m1624 net07701 c32 vss vss nmos L=40e-9 W=90e-9
m1623 net07670 c31 vss vss nmos L=40e-9 W=90e-9
m1622 net07639 c30 vss vss nmos L=40e-9 W=90e-9
m1621 net07608 c29 vss vss nmos L=40e-9 W=90e-9
m1620 net08044 c41 vss vss nmos L=40e-9 W=90e-9
m1619 net08013 net08852 vss vss nmos L=40e-9 W=90e-9
m1618 net07982 c40 vss vss nmos L=40e-9 W=90e-9
m1617 net07951 c39 vss vss nmos L=40e-9 W=90e-9
m1616 net07920 c38 vss vss nmos L=40e-9 W=90e-9
m1615 net07889 c37 vss vss nmos L=40e-9 W=90e-9
m1614 net07858 c36 vss vss nmos L=40e-9 W=90e-9
m1613 net08925 net07826 vss vss nmos L=40e-9 W=90e-9
m1612 net08926 net07795 vss vss nmos L=40e-9 W=90e-9
m1611 net08927 net07764 vss vss nmos L=40e-9 W=90e-9
m1604 net08928 net07733 vss vss nmos L=40e-9 W=90e-9
m1603 net08929 net07702 vss vss nmos L=40e-9 W=90e-9
m1602 net08930 net07671 vss vss nmos L=40e-9 W=90e-9
m1601 net08931 net07640 vss vss nmos L=40e-9 W=90e-9
m1600 net08932 net07609 vss vss nmos L=40e-9 W=90e-9
m1589 net08918 net08045 vss vss nmos L=40e-9 W=90e-9
m1588 net08919 net08014 vss vss nmos L=40e-9 W=90e-9
m1583 net08920 net07983 vss vss nmos L=40e-9 W=90e-9
m1582 net08921 net07952 vss vss nmos L=40e-9 W=90e-9
m1581 net08922 net07921 vss vss nmos L=40e-9 W=90e-9
m1580 net08923 net07890 vss vss nmos L=40e-9 W=90e-9
m1579 net08924 net07859 vss vss nmos L=40e-9 W=90e-9
m1568 net07859 net07832 net08957 vss nmos L=40e-9 W=90e-9
m1567 net07826 net07801 net08958 vss nmos L=40e-9 W=90e-9
m1566 net07795 net07770 net08959 vss nmos L=40e-9 W=90e-9
m1565 net07764 net07739 net08960 vss nmos L=40e-9 W=90e-9
m1564 net07733 net07708 net08961 vss nmos L=40e-9 W=90e-9
m1563 net07702 net07677 net08962 vss nmos L=40e-9 W=90e-9
m1562 net07671 net07646 net08963 vss nmos L=40e-9 W=90e-9
m1561 net07640 net07615 net08964 vss nmos L=40e-9 W=90e-9
m1560 net08076 net08051 net08950 vss nmos L=40e-9 W=90e-9
m1559 net08045 net08020 net08951 vss nmos L=40e-9 W=90e-9
m1558 net08014 net07989 net08952 vss nmos L=40e-9 W=90e-9
m1557 net07983 net07958 net08953 vss nmos L=40e-9 W=90e-9
m1556 net07952 net07927 net08954 vss nmos L=40e-9 W=90e-9
m1555 net07921 net07896 net08955 vss nmos L=40e-9 W=90e-9
m1554 net07890 net07865 net08956 vss nmos L=40e-9 W=90e-9
m1553 net08957 net07834 vss vss nmos L=40e-9 W=90e-9
m1552 net08958 net07803 vss vss nmos L=40e-9 W=90e-9
m1551 net08959 net07772 vss vss nmos L=40e-9 W=90e-9
m1550 net08960 net07741 vss vss nmos L=40e-9 W=90e-9
m1549 net08961 net07710 vss vss nmos L=40e-9 W=90e-9
m1548 net08962 net07679 vss vss nmos L=40e-9 W=90e-9
m1547 net08963 net07648 vss vss nmos L=40e-9 W=90e-9
m1546 net08964 net07617 vss vss nmos L=40e-9 W=90e-9
m1545 net08933 net08584 vss vss nmos L=40e-9 W=90e-9
m1544 net08934 net08553 vss vss nmos L=40e-9 W=90e-9
m1539 net08553 c56 net08966 vss nmos L=40e-9 W=90e-9
m1538 net08584 net08884 net08965 vss nmos L=40e-9 W=90e-9
m1537 net08966 net08528 vss vss nmos L=40e-9 W=90e-9
m1536 net08965 net08559 vss vss nmos L=40e-9 W=90e-9
m1529 net08547 net08541 net09019 vss nmos L=40e-9 W=90e-9
m1528 net08578 net08572 net09017 vss nmos L=40e-9 W=90e-9
m1527 net08572 net08884 vss vss nmos L=40e-9 W=90e-9
m1526 net08541 c56 vss vss nmos L=40e-9 W=90e-9
m1525 net09019 net08528 vss vss nmos L=40e-9 W=90e-9
m1524 net09017 net08559 vss vss nmos L=40e-9 W=90e-9
m1519 net08946 net08179 vss vss nmos L=40e-9 W=90e-9
m1518 net08945 net08210 vss vss nmos L=40e-9 W=90e-9
m1517 net08944 net08241 vss vss nmos L=40e-9 W=90e-9
m1516 net08948 net08117 vss vss nmos L=40e-9 W=90e-9
m1515 net08947 net08148 vss vss nmos L=40e-9 W=90e-9
m1514 net08949 net08084 vss vss nmos L=40e-9 W=90e-9
m1507 net08935 net08522 vss vss nmos L=40e-9 W=90e-9
m1496 net08940 net08367 vss vss nmos L=40e-9 W=90e-9
m1495 net08939 net08398 vss vss nmos L=40e-9 W=90e-9
m1494 net08938 net08429 vss vss nmos L=40e-9 W=90e-9
m1493 net08937 net08460 vss vss nmos L=40e-9 W=90e-9
m1492 net08936 net08491 vss vss nmos L=40e-9 W=90e-9
m1477 net08272 c48 net08975 vss nmos L=40e-9 W=90e-9
m1476 net08303 net08868 net08974 vss nmos L=40e-9 W=90e-9
m1475 net08334 c49 net08973 vss nmos L=40e-9 W=90e-9
m1474 net08117 c43 net08980 vss nmos L=40e-9 W=90e-9
m1473 net08148 c44 net08979 vss nmos L=40e-9 W=90e-9
m1472 net08179 c45 net08978 vss nmos L=40e-9 W=90e-9
m1471 net08210 c46 net08977 vss nmos L=40e-9 W=90e-9
m1470 net08241 c47 net08976 vss nmos L=40e-9 W=90e-9
m1469 net08084 c42 net08981 vss nmos L=40e-9 W=90e-9
m1468 net08522 c55 net08967 vss nmos L=40e-9 W=90e-9
m1467 net08367 c50 net08972 vss nmos L=40e-9 W=90e-9
m1466 net08398 c51 net08971 vss nmos L=40e-9 W=90e-9
m1465 net08429 c52 net08970 vss nmos L=40e-9 W=90e-9
m1464 net08460 c53 net08969 vss nmos L=40e-9 W=90e-9
m1463 net08491 c54 net08968 vss nmos L=40e-9 W=90e-9
m1462 net08975 net08247 vss vss nmos L=40e-9 W=90e-9
m1461 net08974 net08278 vss vss nmos L=40e-9 W=90e-9
m1460 net08973 net08309 vss vss nmos L=40e-9 W=90e-9
m1459 net08980 net08093 vss vss nmos L=40e-9 W=90e-9
m1458 net08979 net08123 vss vss nmos L=40e-9 W=90e-9
m1457 net08978 net08154 vss vss nmos L=40e-9 W=90e-9
m1456 net08977 net08185 vss vss nmos L=40e-9 W=90e-9
m1455 net08976 net08216 vss vss nmos L=40e-9 W=90e-9
m1454 net08981 net08059 vss vss nmos L=40e-9 W=90e-9
m1453 net08967 net08497 vss vss nmos L=40e-9 W=90e-9
m1452 net08972 net08343 vss vss nmos L=40e-9 W=90e-9
m1451 net08971 net08373 vss vss nmos L=40e-9 W=90e-9
m1450 net08970 net08404 vss vss nmos L=40e-9 W=90e-9
m1449 net08969 net08435 vss vss nmos L=40e-9 W=90e-9
m1448 net08968 net08466 vss vss nmos L=40e-9 W=90e-9
m1402 net08266 net08260 net08999 vss nmos L=40e-9 W=90e-9
m1401 net08297 net08291 net08998 vss nmos L=40e-9 W=90e-9
m1400 net08328 net08322 net08997 vss nmos L=40e-9 W=90e-9
m1399 net08111 net08105 net09004 vss nmos L=40e-9 W=90e-9
m1398 net08142 net08136 net09003 vss nmos L=40e-9 W=90e-9
m1397 net08173 net08167 net09002 vss nmos L=40e-9 W=90e-9
m1396 net08204 net08198 net09001 vss nmos L=40e-9 W=90e-9
m1395 net08235 net08229 net09000 vss nmos L=40e-9 W=90e-9
m1394 net08078 net08072 net09005 vss nmos L=40e-9 W=90e-9
m1393 net08516 net08510 net09021 vss nmos L=40e-9 W=90e-9
m1392 net08485 net08479 net09023 vss nmos L=40e-9 W=90e-9
m1391 net08454 net08448 net09025 vss nmos L=40e-9 W=90e-9
m1390 net08423 net08417 net09027 vss nmos L=40e-9 W=90e-9
m1389 net08392 net08386 net09029 vss nmos L=40e-9 W=90e-9
m1388 net08361 net08355 net09031 vss nmos L=40e-9 W=90e-9
m1387 net08260 c48 vss vss nmos L=40e-9 W=90e-9
m1386 net08291 net08868 vss vss nmos L=40e-9 W=90e-9
m1385 net08322 c49 vss vss nmos L=40e-9 W=90e-9
m1384 net08105 c43 vss vss nmos L=40e-9 W=90e-9
m1383 net08136 c44 vss vss nmos L=40e-9 W=90e-9
m1382 net08167 c45 vss vss nmos L=40e-9 W=90e-9
m1381 net08198 c46 vss vss nmos L=40e-9 W=90e-9
m1380 net08229 c47 vss vss nmos L=40e-9 W=90e-9
m1379 net08072 c42 vss vss nmos L=40e-9 W=90e-9
m1378 net08510 c55 vss vss nmos L=40e-9 W=90e-9
m1377 net08479 c54 vss vss nmos L=40e-9 W=90e-9
m1376 net08448 c53 vss vss nmos L=40e-9 W=90e-9
m1375 net08417 c52 vss vss nmos L=40e-9 W=90e-9
m1374 net08386 c51 vss vss nmos L=40e-9 W=90e-9
m1373 net08355 c50 vss vss nmos L=40e-9 W=90e-9
m1372 net08999 net08247 vss vss nmos L=40e-9 W=90e-9
m1371 net08998 net08278 vss vss nmos L=40e-9 W=90e-9
m1370 net08997 net08309 vss vss nmos L=40e-9 W=90e-9
m1369 net09004 net08093 vss vss nmos L=40e-9 W=90e-9
m1368 net09003 net08123 vss vss nmos L=40e-9 W=90e-9
m1367 net09002 net08154 vss vss nmos L=40e-9 W=90e-9
m1366 net09001 net08185 vss vss nmos L=40e-9 W=90e-9
m1365 net09000 net08216 vss vss nmos L=40e-9 W=90e-9
m1358 net09005 net08059 vss vss nmos L=40e-9 W=90e-9
m1345 net09021 net08497 vss vss nmos L=40e-9 W=90e-9
m1342 net09023 net08466 vss vss nmos L=40e-9 W=90e-9
m1341 net09025 net08435 vss vss nmos L=40e-9 W=90e-9
m1340 net09027 net08404 vss vss nmos L=40e-9 W=90e-9
m1339 net09029 net08373 vss vss nmos L=40e-9 W=90e-9
m1338 net09031 net08343 vss vss nmos L=40e-9 W=90e-9
m1327 net08950 net08053 vss vss nmos L=40e-9 W=90e-9
m1326 net08951 net08022 vss vss nmos L=40e-9 W=90e-9
m1319 net08952 net07991 vss vss nmos L=40e-9 W=90e-9
m1318 net08953 net07960 vss vss nmos L=40e-9 W=90e-9
m1317 net08954 net07929 vss vss nmos L=40e-9 W=90e-9
m1316 net08955 net07898 vss vss nmos L=40e-9 W=90e-9
m1315 net08956 net07867 vss vss nmos L=40e-9 W=90e-9
m1290 net07834 c35 net08989 vss nmos L=40e-9 W=90e-9
m1289 net07803 c34 net08990 vss nmos L=40e-9 W=90e-9
m1288 net07772 c33 net08991 vss nmos L=40e-9 W=90e-9
m1287 net07741 net08836 net08992 vss nmos L=40e-9 W=90e-9
m1286 net07710 c32 net08993 vss nmos L=40e-9 W=90e-9
m1285 net07679 c31 net08994 vss nmos L=40e-9 W=90e-9
m1284 net07648 c30 net08995 vss nmos L=40e-9 W=90e-9
m1283 net07617 c29 net08996 vss nmos L=40e-9 W=90e-9
m1282 net08053 c41 net08982 vss nmos L=40e-9 W=90e-9
m1281 net08022 net08852 net08983 vss nmos L=40e-9 W=90e-9
m1280 net07991 c40 net08984 vss nmos L=40e-9 W=90e-9
m1279 net07960 c39 net08985 vss nmos L=40e-9 W=90e-9
m1278 net07929 c38 net08986 vss nmos L=40e-9 W=90e-9
m1277 net07898 c37 net08987 vss nmos L=40e-9 W=90e-9
m1276 net07867 c36 net08988 vss nmos L=40e-9 W=90e-9
m1275 net08989 net07809 vss vss nmos L=40e-9 W=90e-9
m1274 net08990 net07778 vss vss nmos L=40e-9 W=90e-9
m1273 net08991 net07747 vss vss nmos L=40e-9 W=90e-9
m1272 net08992 net07716 vss vss nmos L=40e-9 W=90e-9
m1271 net08993 net07685 vss vss nmos L=40e-9 W=90e-9
m1270 net08994 net07654 vss vss nmos L=40e-9 W=90e-9
m1269 net08995 net07623 vss vss nmos L=40e-9 W=90e-9
m1268 net08996 net07593 vss vss nmos L=40e-9 W=90e-9
m1267 net08982 net08028 vss vss nmos L=40e-9 W=90e-9
m1266 net08983 net07997 vss vss nmos L=40e-9 W=90e-9
m1265 net08984 net07966 vss vss nmos L=40e-9 W=90e-9
m1264 net08985 net07935 vss vss nmos L=40e-9 W=90e-9
m1263 net08986 net07904 vss vss nmos L=40e-9 W=90e-9
m1262 net08987 net07873 vss vss nmos L=40e-9 W=90e-9
m1261 net08988 net07843 vss vss nmos L=40e-9 W=90e-9
m1215 net07828 net07822 net09008 vss nmos L=40e-9 W=90e-9
m1214 net07797 net07791 net09009 vss nmos L=40e-9 W=90e-9
m1213 net07766 net07760 net09010 vss nmos L=40e-9 W=90e-9
m1212 net07735 net07729 net09011 vss nmos L=40e-9 W=90e-9
m1211 net07704 net07698 net09012 vss nmos L=40e-9 W=90e-9
m1210 net07673 net07667 net09013 vss nmos L=40e-9 W=90e-9
m1209 net07642 net07636 net09014 vss nmos L=40e-9 W=90e-9
m1208 net07611 net07605 net09015 vss nmos L=40e-9 W=90e-9
m1207 net08016 net08010 net09007 vss nmos L=40e-9 W=90e-9
m1206 net08047 net08041 net09006 vss nmos L=40e-9 W=90e-9
m1205 net07861 net07855 net09052 vss nmos L=40e-9 W=90e-9
m1204 net07892 net07886 net09050 vss nmos L=40e-9 W=90e-9
m1203 net07923 net07917 net09048 vss nmos L=40e-9 W=90e-9
m1202 net07954 net07948 net09046 vss nmos L=40e-9 W=90e-9
m1201 net07985 net07979 net09044 vss nmos L=40e-9 W=90e-9
m1200 net07822 c35 vss vss nmos L=40e-9 W=90e-9
m1199 net07791 c34 vss vss nmos L=40e-9 W=90e-9
m1198 net07760 c33 vss vss nmos L=40e-9 W=90e-9
m1197 net07729 net08836 vss vss nmos L=40e-9 W=90e-9
m1196 net07698 c32 vss vss nmos L=40e-9 W=90e-9
m1195 net07667 c31 vss vss nmos L=40e-9 W=90e-9
m1194 net07636 c30 vss vss nmos L=40e-9 W=90e-9
m1193 net07605 c29 vss vss nmos L=40e-9 W=90e-9
m1192 net08010 net08852 vss vss nmos L=40e-9 W=90e-9
m1191 net08041 c41 vss vss nmos L=40e-9 W=90e-9
m1190 net07855 c36 vss vss nmos L=40e-9 W=90e-9
m1189 net07886 c37 vss vss nmos L=40e-9 W=90e-9
m1188 net07917 c38 vss vss nmos L=40e-9 W=90e-9
m1187 net07948 c39 vss vss nmos L=40e-9 W=90e-9
m1186 net07979 c40 vss vss nmos L=40e-9 W=90e-9
m1185 net09008 net07809 vss vss nmos L=40e-9 W=90e-9
m1184 net09009 net07778 vss vss nmos L=40e-9 W=90e-9
m1183 net09010 net07747 vss vss nmos L=40e-9 W=90e-9
m1176 net09011 net07716 vss vss nmos L=40e-9 W=90e-9
m1175 net09012 net07685 vss vss nmos L=40e-9 W=90e-9
m1174 net09013 net07654 vss vss nmos L=40e-9 W=90e-9
m1173 net09014 net07623 vss vss nmos L=40e-9 W=90e-9
m1172 net09015 net07593 vss vss nmos L=40e-9 W=90e-9
m1161 net09007 net07997 vss vss nmos L=40e-9 W=90e-9
m1160 net09006 net08028 vss vss nmos L=40e-9 W=90e-9
m1159 net09052 net07843 vss vss nmos L=40e-9 W=90e-9
m1158 net09050 net07873 vss vss nmos L=40e-9 W=90e-9
m1157 net09048 net07904 vss vss nmos L=40e-9 W=90e-9
m1156 net09046 net07935 vss vss nmos L=40e-9 W=90e-9
m1155 net09044 net07966 vss vss nmos L=40e-9 W=90e-9
m1140 net08593 net08578 net09016 vss nmos L=40e-9 W=90e-9
m1139 net08559 net08547 net09018 vss nmos L=40e-9 W=90e-9
m1138 net09018 net08549 vss vss nmos L=40e-9 W=90e-9
m1137 net09016 net08580 vss vss nmos L=40e-9 W=90e-9
m1132 net08549 c56 net09062 vss nmos L=40e-9 W=90e-9
m1131 net08580 net08884 net09061 vss nmos L=40e-9 W=90e-9
m1130 net09062 net08545 vss vss nmos L=40e-9 W=90e-9
m1129 net09061 net08576 vss vss nmos L=40e-9 W=90e-9
m1128 net08309 net08297 net09033 vss nmos L=40e-9 W=90e-9
m1127 net08343 net08328 net09032 vss nmos L=40e-9 W=90e-9
m1126 net08278 net08266 net09034 vss nmos L=40e-9 W=90e-9
m1125 net08123 net08111 net09039 vss nmos L=40e-9 W=90e-9
m1124 net08154 net08142 net09038 vss nmos L=40e-9 W=90e-9
m1123 net08185 net08173 net09037 vss nmos L=40e-9 W=90e-9
m1122 net08216 net08204 net09036 vss nmos L=40e-9 W=90e-9
m1121 net08247 net08235 net09035 vss nmos L=40e-9 W=90e-9
m1120 net08093 net08078 net09040 vss nmos L=40e-9 W=90e-9
m1119 net08528 net08516 net09020 vss nmos L=40e-9 W=90e-9
m1118 net08497 net08485 net09022 vss nmos L=40e-9 W=90e-9
m1117 net08466 net08454 net09024 vss nmos L=40e-9 W=90e-9
m1116 net08435 net08423 net09026 vss nmos L=40e-9 W=90e-9
m1115 net08404 net08392 net09028 vss nmos L=40e-9 W=90e-9
m1114 net08373 net08361 net09030 vss nmos L=40e-9 W=90e-9
m1113 net09034 net08268 vss vss nmos L=40e-9 W=90e-9
m1112 net09033 net08299 vss vss nmos L=40e-9 W=90e-9
m1111 net09032 net08330 vss vss nmos L=40e-9 W=90e-9
m1110 net09039 net08113 vss vss nmos L=40e-9 W=90e-9
m1109 net09038 net08144 vss vss nmos L=40e-9 W=90e-9
m1108 net09037 net08175 vss vss nmos L=40e-9 W=90e-9
m1107 net09036 net08206 vss vss nmos L=40e-9 W=90e-9
m1106 net09035 net08237 vss vss nmos L=40e-9 W=90e-9
m1105 net09040 net08080 vss vss nmos L=40e-9 W=90e-9
m1098 net09020 net08518 vss vss nmos L=40e-9 W=90e-9
m1087 net09022 net08487 vss vss nmos L=40e-9 W=90e-9
m1086 net09024 net08456 vss vss nmos L=40e-9 W=90e-9
m1085 net09026 net08425 vss vss nmos L=40e-9 W=90e-9
m1084 net09028 net08394 vss vss nmos L=40e-9 W=90e-9
m1083 net09030 net08363 vss vss nmos L=40e-9 W=90e-9
m1068 net08268 c48 net09071 vss nmos L=40e-9 W=90e-9
m1067 net08299 net08868 net09070 vss nmos L=40e-9 W=90e-9
m1066 net08330 c49 net09069 vss nmos L=40e-9 W=90e-9
m1065 net08113 c43 net09076 vss nmos L=40e-9 W=90e-9
m1064 net08144 c44 net09075 vss nmos L=40e-9 W=90e-9
m1063 net08175 c45 net09074 vss nmos L=40e-9 W=90e-9
m1062 net08206 c46 net09073 vss nmos L=40e-9 W=90e-9
m1061 net08237 c47 net09072 vss nmos L=40e-9 W=90e-9
m1060 net08080 c42 net09077 vss nmos L=40e-9 W=90e-9
m1059 net08518 c55 net09063 vss nmos L=40e-9 W=90e-9
m1058 net08487 c54 net09064 vss nmos L=40e-9 W=90e-9
m1057 net08456 c53 net09065 vss nmos L=40e-9 W=90e-9
m1056 net08425 c52 net09066 vss nmos L=40e-9 W=90e-9
m1055 net08394 c51 net09067 vss nmos L=40e-9 W=90e-9
m1054 net08363 c50 net09068 vss nmos L=40e-9 W=90e-9
m1053 net09071 net08264 vss vss nmos L=40e-9 W=90e-9
m1052 net09070 net08295 vss vss nmos L=40e-9 W=90e-9
m1051 net09069 net08326 vss vss nmos L=40e-9 W=90e-9
m1050 net09076 net08109 vss vss nmos L=40e-9 W=90e-9
m1049 net09075 net08140 vss vss nmos L=40e-9 W=90e-9
m1048 net09074 net08171 vss vss nmos L=40e-9 W=90e-9
m1047 net09073 net08202 vss vss nmos L=40e-9 W=90e-9
m1046 net09072 net08233 vss vss nmos L=40e-9 W=90e-9
m1045 net09077 net08076 vss vss nmos L=40e-9 W=90e-9
m1044 net09063 net08514 vss vss nmos L=40e-9 W=90e-9
m1043 net09068 net08359 vss vss nmos L=40e-9 W=90e-9
m1042 net09064 net08483 vss vss nmos L=40e-9 W=90e-9
m1041 net09065 net08452 vss vss nmos L=40e-9 W=90e-9
m1040 net09066 net08421 vss vss nmos L=40e-9 W=90e-9
m1039 net09067 net08390 vss vss nmos L=40e-9 W=90e-9
m1038 net07843 net07828 net09053 vss nmos L=40e-9 W=90e-9
m1037 net07809 net07797 net09054 vss nmos L=40e-9 W=90e-9
m1036 net07778 net07766 net09055 vss nmos L=40e-9 W=90e-9
m1035 net07747 net07735 net09056 vss nmos L=40e-9 W=90e-9
m1034 net07716 net07704 net09057 vss nmos L=40e-9 W=90e-9
m1033 net07685 net07673 net09058 vss nmos L=40e-9 W=90e-9
m1032 net07654 net07642 net09059 vss nmos L=40e-9 W=90e-9
m1031 net07623 net07611 net09060 vss nmos L=40e-9 W=90e-9
m1030 net08028 net08016 net09042 vss nmos L=40e-9 W=90e-9
m1029 net08059 net08047 net09041 vss nmos L=40e-9 W=90e-9
m1028 net07873 net07861 net09051 vss nmos L=40e-9 W=90e-9
m1027 net07904 net07892 net09049 vss nmos L=40e-9 W=90e-9
m1026 net07935 net07923 net09047 vss nmos L=40e-9 W=90e-9
m1025 net07966 net07954 net09045 vss nmos L=40e-9 W=90e-9
m1024 net07997 net07985 net09043 vss nmos L=40e-9 W=90e-9
m1023 net09053 net07830 vss vss nmos L=40e-9 W=90e-9
m1022 net09054 net07799 vss vss nmos L=40e-9 W=90e-9
m1021 net09055 net07768 vss vss nmos L=40e-9 W=90e-9
m1020 net09056 net07737 vss vss nmos L=40e-9 W=90e-9
m1019 net09057 net07706 vss vss nmos L=40e-9 W=90e-9
m1018 net09058 net07675 vss vss nmos L=40e-9 W=90e-9
m1017 net09059 net07644 vss vss nmos L=40e-9 W=90e-9
m1016 net09060 net07613 vss vss nmos L=40e-9 W=90e-9
m1015 net09042 net08018 vss vss nmos L=40e-9 W=90e-9
m1014 net09041 net08049 vss vss nmos L=40e-9 W=90e-9
m1007 net09051 net07863 vss vss nmos L=40e-9 W=90e-9
m1006 net09049 net07894 vss vss nmos L=40e-9 W=90e-9
m1005 net09047 net07925 vss vss nmos L=40e-9 W=90e-9
m1004 net09045 net07956 vss vss nmos L=40e-9 W=90e-9
m1003 net09043 net07987 vss vss nmos L=40e-9 W=90e-9
m978 net07830 c35 net09085 vss nmos L=40e-9 W=90e-9
m977 net07799 c34 net09086 vss nmos L=40e-9 W=90e-9
m976 net07768 c33 net09087 vss nmos L=40e-9 W=90e-9
m975 net07737 net08836 net09088 vss nmos L=40e-9 W=90e-9
m974 net07706 c32 net09089 vss nmos L=40e-9 W=90e-9
m973 net07675 c31 net09090 vss nmos L=40e-9 W=90e-9
m972 net07644 c30 net09091 vss nmos L=40e-9 W=90e-9
m971 net07613 c29 net09092 vss nmos L=40e-9 W=90e-9
m970 net08018 net08852 net09079 vss nmos L=40e-9 W=90e-9
m969 net08049 c41 net09078 vss nmos L=40e-9 W=90e-9
m968 net07863 c36 net09084 vss nmos L=40e-9 W=90e-9
m967 net07894 c37 net09083 vss nmos L=40e-9 W=90e-9
m966 net07925 c38 net09082 vss nmos L=40e-9 W=90e-9
m965 net07956 c39 net09081 vss nmos L=40e-9 W=90e-9
m964 net07987 c40 net09080 vss nmos L=40e-9 W=90e-9
m963 net09085 net07826 vss vss nmos L=40e-9 W=90e-9
m962 net09086 net07795 vss vss nmos L=40e-9 W=90e-9
m961 net09087 net07764 vss vss nmos L=40e-9 W=90e-9
m960 net09088 net07733 vss vss nmos L=40e-9 W=90e-9
m959 net09089 net07702 vss vss nmos L=40e-9 W=90e-9
m958 net09090 net07671 vss vss nmos L=40e-9 W=90e-9
m957 net09091 net07640 vss vss nmos L=40e-9 W=90e-9
m956 net09092 net07609 vss vss nmos L=40e-9 W=90e-9
m955 net09079 net08014 vss vss nmos L=40e-9 W=90e-9
m954 net09078 net08045 vss vss nmos L=40e-9 W=90e-9
m953 net09083 net07890 vss vss nmos L=40e-9 W=90e-9
m952 net09082 net07921 vss vss nmos L=40e-9 W=90e-9
m951 net09081 net07952 vss vss nmos L=40e-9 W=90e-9
m950 net09080 net07983 vss vss nmos L=40e-9 W=90e-9
m949 net09084 net07859 vss vss nmos L=40e-9 W=90e-9
m947 net09109 net07584 vss vss nmos L=40e-9 W=90e-9
m946 net07609 net07582 net09109 vss nmos L=40e-9 W=90e-9
m942 net07584 c28 net09110 vss nmos L=40e-9 W=90e-9
m941 net09110 net07559 vss vss nmos L=40e-9 W=90e-9
m940 net09093 net07576 vss vss nmos L=40e-9 W=90e-9
m939 net07582 net07575 net09093 vss nmos L=40e-9 W=90e-9
m936 net07575 c28 vss vss nmos L=40e-9 W=90e-9
m933 net09111 net07552 vss vss nmos L=40e-9 W=90e-9
m932 net07576 net07550 net09111 vss nmos L=40e-9 W=90e-9
m928 net09112 net07527 vss vss nmos L=40e-9 W=90e-9
m927 net07552 c27 net09112 vss nmos L=40e-9 W=90e-9
m926 net09094 net07544 vss vss nmos L=40e-9 W=90e-9
m925 net07550 net07543 net09094 vss nmos L=40e-9 W=90e-9
m922 net07543 c27 vss vss nmos L=40e-9 W=90e-9
m919 net09113 net07520 vss vss nmos L=40e-9 W=90e-9
m918 net07544 net07518 net09113 vss nmos L=40e-9 W=90e-9
m914 net09114 net07494 vss vss nmos L=40e-9 W=90e-9
m913 net07520 c26 net09114 vss nmos L=40e-9 W=90e-9
m912 net09095 net07511 vss vss nmos L=40e-9 W=90e-9
m911 net07518 net07510 net09095 vss nmos L=40e-9 W=90e-9
m908 net07510 c26 vss vss nmos L=40e-9 W=90e-9
m905 net09115 net07488 vss vss nmos L=40e-9 W=90e-9
m904 net07511 net07486 net09115 vss nmos L=40e-9 W=90e-9
m900 net09116 net07463 vss vss nmos L=40e-9 W=90e-9
m899 net07488 c25 net09116 vss nmos L=40e-9 W=90e-9
m898 net09096 net07480 vss vss nmos L=40e-9 W=90e-9
m897 net07486 net07479 net09096 vss nmos L=40e-9 W=90e-9
m894 net07479 c25 vss vss nmos L=40e-9 W=90e-9
m891 net09117 net07457 vss vss nmos L=40e-9 W=90e-9
m890 net07480 net07455 net09117 vss nmos L=40e-9 W=90e-9
m886 net09118 net07432 vss vss nmos L=40e-9 W=90e-9
m885 net07457 net08819 net09118 vss nmos L=40e-9 W=90e-9
m884 net09097 net07449 vss vss nmos L=40e-9 W=90e-9
m883 net07455 net07448 net09097 vss nmos L=40e-9 W=90e-9
m880 net07448 net08819 vss vss nmos L=40e-9 W=90e-9
m877 net09119 net07426 vss vss nmos L=40e-9 W=90e-9
m876 net07449 net07424 net09119 vss nmos L=40e-9 W=90e-9
m872 net09120 net07401 vss vss nmos L=40e-9 W=90e-9
m871 net07426 c24 net09120 vss nmos L=40e-9 W=90e-9
m870 net09098 net07418 vss vss nmos L=40e-9 W=90e-9
m869 net07424 net07417 net09098 vss nmos L=40e-9 W=90e-9
m866 net07417 c24 vss vss nmos L=40e-9 W=90e-9
m863 net09121 net07395 vss vss nmos L=40e-9 W=90e-9
m862 net07418 net07393 net09121 vss nmos L=40e-9 W=90e-9
m858 net09122 net07370 vss vss nmos L=40e-9 W=90e-9
m857 net07395 c23 net09122 vss nmos L=40e-9 W=90e-9
m856 net09099 net07387 vss vss nmos L=40e-9 W=90e-9
m855 net07393 net07386 net09099 vss nmos L=40e-9 W=90e-9
m852 net07386 c23 vss vss nmos L=40e-9 W=90e-9
m849 net09123 net07364 vss vss nmos L=40e-9 W=90e-9
m848 net07387 net07362 net09123 vss nmos L=40e-9 W=90e-9
m844 net07364 c22 net09124 vss nmos L=40e-9 W=90e-9
m843 net09124 net07340 vss vss nmos L=40e-9 W=90e-9
m842 net09100 net07356 vss vss nmos L=40e-9 W=90e-9
m841 net07362 net07355 net09100 vss nmos L=40e-9 W=90e-9
m838 net07355 c22 vss vss nmos L=40e-9 W=90e-9
m812 net07329 net07322 net09101 vss nmos L=40e-9 W=90e-9
m811 net07298 net07291 net09102 vss nmos L=40e-9 W=90e-9
m810 net07267 net07260 net09103 vss nmos L=40e-9 W=90e-9
m809 net07236 net07228 net09104 vss nmos L=40e-9 W=90e-9
m808 net07204 net07197 net09105 vss nmos L=40e-9 W=90e-9
m807 net07173 net07166 net09106 vss nmos L=40e-9 W=90e-9
m806 net07142 net07135 net09107 vss nmos L=40e-9 W=90e-9
m805 net07111 net07104 net09108 vss nmos L=40e-9 W=90e-9
m804 net07322 c21 vss vss nmos L=40e-9 W=90e-9
m803 net07291 c20 vss vss nmos L=40e-9 W=90e-9
m802 net07260 c19 vss vss nmos L=40e-9 W=90e-9
m801 net07228 c18 vss vss nmos L=40e-9 W=90e-9
m800 net07197 c17 vss vss nmos L=40e-9 W=90e-9
m799 net07166 net08803 vss vss nmos L=40e-9 W=90e-9
m798 net07135 c16 vss vss nmos L=40e-9 W=90e-9
m797 net07104 c15 vss vss nmos L=40e-9 W=90e-9
m796 net09101 net07323 vss vss nmos L=40e-9 W=90e-9
m795 net09102 net07292 vss vss nmos L=40e-9 W=90e-9
m794 net09103 net07261 vss vss nmos L=40e-9 W=90e-9
m787 net09104 net07229 vss vss nmos L=40e-9 W=90e-9
m786 net09105 net07198 vss vss nmos L=40e-9 W=90e-9
m785 net09106 net07167 vss vss nmos L=40e-9 W=90e-9
m784 net09107 net07136 vss vss nmos L=40e-9 W=90e-9
m783 net09108 net07105 vss vss nmos L=40e-9 W=90e-9
m772 net07356 net07329 net09125 vss nmos L=40e-9 W=90e-9
m771 net07323 net07298 net09127 vss nmos L=40e-9 W=90e-9
m770 net07292 net07267 net09129 vss nmos L=40e-9 W=90e-9
m769 net07261 net07236 net09131 vss nmos L=40e-9 W=90e-9
m768 net07229 net07204 net09133 vss nmos L=40e-9 W=90e-9
m767 net07198 net07173 net09135 vss nmos L=40e-9 W=90e-9
m766 net07167 net07142 net09137 vss nmos L=40e-9 W=90e-9
m765 net07136 net07111 net09139 vss nmos L=40e-9 W=90e-9
m764 net09125 net07331 vss vss nmos L=40e-9 W=90e-9
m763 net09127 net07300 vss vss nmos L=40e-9 W=90e-9
m762 net09129 net07269 vss vss nmos L=40e-9 W=90e-9
m761 net09131 net07238 vss vss nmos L=40e-9 W=90e-9
m760 net09133 net07206 vss vss nmos L=40e-9 W=90e-9
m759 net09135 net07175 vss vss nmos L=40e-9 W=90e-9
m758 net09137 net07144 vss vss nmos L=40e-9 W=90e-9
m757 net09139 net07113 vss vss nmos L=40e-9 W=90e-9
m740 net07331 c21 net09126 vss nmos L=40e-9 W=90e-9
m739 net07300 c20 net09128 vss nmos L=40e-9 W=90e-9
m738 net07269 c19 net09130 vss nmos L=40e-9 W=90e-9
m737 net07238 c18 net09132 vss nmos L=40e-9 W=90e-9
m736 net07206 c17 net09134 vss nmos L=40e-9 W=90e-9
m735 net07175 net08803 net09136 vss nmos L=40e-9 W=90e-9
m734 net07144 c16 net09138 vss nmos L=40e-9 W=90e-9
m733 net07113 c15 net09140 vss nmos L=40e-9 W=90e-9
m732 net09126 net07306 vss vss nmos L=40e-9 W=90e-9
m731 net09128 net07275 vss vss nmos L=40e-9 W=90e-9
m730 net09130 net07244 vss vss nmos L=40e-9 W=90e-9
m729 net09132 net07212 vss vss nmos L=40e-9 W=90e-9
m728 net09134 net07181 vss vss nmos L=40e-9 W=90e-9
m727 net09136 net07150 vss vss nmos L=40e-9 W=90e-9
m726 net09138 net07119 vss vss nmos L=40e-9 W=90e-9
m725 net09140 net07089 vss vss nmos L=40e-9 W=90e-9
m722 net07578 net07572 net09142 vss nmos L=40e-9 W=90e-9
m721 net09142 net07559 vss vss nmos L=40e-9 W=90e-9
m718 net07593 net07578 net09141 vss nmos L=40e-9 W=90e-9
m717 net09141 net07580 vss vss nmos L=40e-9 W=90e-9
m714 net07580 c28 net09173 vss nmos L=40e-9 W=90e-9
m713 net09173 net07576 vss vss nmos L=40e-9 W=90e-9
m690 net07513 net07507 net09146 vss nmos L=40e-9 W=90e-9
m689 net07546 net07540 net09144 vss nmos L=40e-9 W=90e-9
m688 net07358 net07352 net09156 vss nmos L=40e-9 W=90e-9
m687 net07389 net07383 net09154 vss nmos L=40e-9 W=90e-9
m686 net07420 net07414 net09152 vss nmos L=40e-9 W=90e-9
m685 net07451 net07445 net09150 vss nmos L=40e-9 W=90e-9
m684 net07482 net07476 net09148 vss nmos L=40e-9 W=90e-9
m683 net07507 c26 vss vss nmos L=40e-9 W=90e-9
m682 net07540 c27 vss vss nmos L=40e-9 W=90e-9
m681 net07572 c28 vss vss nmos L=40e-9 W=90e-9
m680 net07352 c22 vss vss nmos L=40e-9 W=90e-9
m679 net07383 c23 vss vss nmos L=40e-9 W=90e-9
m678 net07414 c24 vss vss nmos L=40e-9 W=90e-9
m677 net07445 net08819 vss vss nmos L=40e-9 W=90e-9
m676 net07476 c25 vss vss nmos L=40e-9 W=90e-9
m675 net09146 net07494 vss vss nmos L=40e-9 W=90e-9
m674 net09144 net07527 vss vss nmos L=40e-9 W=90e-9
m673 net09156 net07340 vss vss nmos L=40e-9 W=90e-9
m672 net09154 net07370 vss vss nmos L=40e-9 W=90e-9
m671 net09152 net07401 vss vss nmos L=40e-9 W=90e-9
m670 net09150 net07432 vss vss nmos L=40e-9 W=90e-9
m669 net09148 net07463 vss vss nmos L=40e-9 W=90e-9
m654 net07527 net07513 net09145 vss nmos L=40e-9 W=90e-9
m653 net07559 net07546 net09143 vss nmos L=40e-9 W=90e-9
m652 net07370 net07358 net09155 vss nmos L=40e-9 W=90e-9
m651 net07401 net07389 net09153 vss nmos L=40e-9 W=90e-9
m650 net07432 net07420 net09151 vss nmos L=40e-9 W=90e-9
m649 net07463 net07451 net09149 vss nmos L=40e-9 W=90e-9
m648 net07494 net07482 net09147 vss nmos L=40e-9 W=90e-9
m647 net09145 net07516 vss vss nmos L=40e-9 W=90e-9
m646 net09143 net07548 vss vss nmos L=40e-9 W=90e-9
m645 net09155 net07360 vss vss nmos L=40e-9 W=90e-9
m644 net09153 net07391 vss vss nmos L=40e-9 W=90e-9
m643 net09151 net07422 vss vss nmos L=40e-9 W=90e-9
m642 net09149 net07453 vss vss nmos L=40e-9 W=90e-9
m641 net09147 net07484 vss vss nmos L=40e-9 W=90e-9
m626 net07516 c26 net09175 vss nmos L=40e-9 W=90e-9
m625 net07548 c27 net09174 vss nmos L=40e-9 W=90e-9
m624 net07360 c22 net09180 vss nmos L=40e-9 W=90e-9
m623 net07391 c23 net09179 vss nmos L=40e-9 W=90e-9
m622 net07422 c24 net09178 vss nmos L=40e-9 W=90e-9
m621 net07453 net08819 net09177 vss nmos L=40e-9 W=90e-9
m620 net07484 c25 net09176 vss nmos L=40e-9 W=90e-9
m619 net09175 net07511 vss vss nmos L=40e-9 W=90e-9
m618 net09174 net07544 vss vss nmos L=40e-9 W=90e-9
m617 net09179 net07387 vss vss nmos L=40e-9 W=90e-9
m616 net09178 net07418 vss vss nmos L=40e-9 W=90e-9
m615 net09177 net07449 vss vss nmos L=40e-9 W=90e-9
m614 net09176 net07480 vss vss nmos L=40e-9 W=90e-9
m613 net09180 net07356 vss vss nmos L=40e-9 W=90e-9
m588 net07325 net07319 net09158 vss nmos L=40e-9 W=90e-9
m587 net07294 net07288 net09160 vss nmos L=40e-9 W=90e-9
m586 net07263 net07257 net09162 vss nmos L=40e-9 W=90e-9
m585 net07231 net07225 net09164 vss nmos L=40e-9 W=90e-9
m584 net07200 net07194 net09166 vss nmos L=40e-9 W=90e-9
m583 net07169 net07163 net09168 vss nmos L=40e-9 W=90e-9
m582 net07138 net07132 net09170 vss nmos L=40e-9 W=90e-9
m581 net07107 net07101 net09172 vss nmos L=40e-9 W=90e-9
m580 net07319 c21 vss vss nmos L=40e-9 W=90e-9
m579 net07288 c20 vss vss nmos L=40e-9 W=90e-9
m578 net07257 c19 vss vss nmos L=40e-9 W=90e-9
m577 net07225 c18 vss vss nmos L=40e-9 W=90e-9
m576 net07194 c17 vss vss nmos L=40e-9 W=90e-9
m575 net07163 net08803 vss vss nmos L=40e-9 W=90e-9
m574 net07132 c16 vss vss nmos L=40e-9 W=90e-9
m573 net07101 c15 vss vss nmos L=40e-9 W=90e-9
m572 net09158 net07306 vss vss nmos L=40e-9 W=90e-9
m571 net09160 net07275 vss vss nmos L=40e-9 W=90e-9
m570 net09162 net07244 vss vss nmos L=40e-9 W=90e-9
m563 net09164 net07212 vss vss nmos L=40e-9 W=90e-9
m562 net09166 net07181 vss vss nmos L=40e-9 W=90e-9
m561 net09168 net07150 vss vss nmos L=40e-9 W=90e-9
m560 net09170 net07119 vss vss nmos L=40e-9 W=90e-9
m559 net09172 net07089 vss vss nmos L=40e-9 W=90e-9
m548 net07340 net07325 net09157 vss nmos L=40e-9 W=90e-9
m547 net07306 net07294 net09159 vss nmos L=40e-9 W=90e-9
m546 net07275 net07263 net09161 vss nmos L=40e-9 W=90e-9
m545 net07244 net07231 net09163 vss nmos L=40e-9 W=90e-9
m544 net07212 net07200 net09165 vss nmos L=40e-9 W=90e-9
m543 net07181 net07169 net09167 vss nmos L=40e-9 W=90e-9
m542 net07150 net07138 net09169 vss nmos L=40e-9 W=90e-9
m541 net07119 net07107 net09171 vss nmos L=40e-9 W=90e-9
m540 net09157 net07327 vss vss nmos L=40e-9 W=90e-9
m539 net09159 net07296 vss vss nmos L=40e-9 W=90e-9
m538 net09161 net07265 vss vss nmos L=40e-9 W=90e-9
m537 net09163 net07234 vss vss nmos L=40e-9 W=90e-9
m536 net09165 net07202 vss vss nmos L=40e-9 W=90e-9
m535 net09167 net07171 vss vss nmos L=40e-9 W=90e-9
m534 net09169 net07140 vss vss nmos L=40e-9 W=90e-9
m533 net09171 net07109 vss vss nmos L=40e-9 W=90e-9
m516 net07327 c21 net09181 vss nmos L=40e-9 W=90e-9
m515 net07296 c20 net09182 vss nmos L=40e-9 W=90e-9
m514 net07265 c19 net09183 vss nmos L=40e-9 W=90e-9
m513 net07234 c18 net09184 vss nmos L=40e-9 W=90e-9
m512 net07202 c17 net09185 vss nmos L=40e-9 W=90e-9
m511 net07171 net08803 net09186 vss nmos L=40e-9 W=90e-9
m510 net07140 c16 net09187 vss nmos L=40e-9 W=90e-9
m509 net07109 c15 net09188 vss nmos L=40e-9 W=90e-9
m508 net09181 net07323 vss vss nmos L=40e-9 W=90e-9
m507 net09182 net07292 vss vss nmos L=40e-9 W=90e-9
m506 net09183 net07261 vss vss nmos L=40e-9 W=90e-9
m505 net09184 net07229 vss vss nmos L=40e-9 W=90e-9
m504 net09185 net07198 vss vss nmos L=40e-9 W=90e-9
m503 net09186 net07167 vss vss nmos L=40e-9 W=90e-9
m502 net09187 net07136 vss vss nmos L=40e-9 W=90e-9
m501 net09188 net07105 vss vss nmos L=40e-9 W=90e-9
m492 net07076 net07067 net09190 vss nmos L=40e-9 W=90e-9
m491 net07041 net07033 net09192 vss nmos L=40e-9 W=90e-9
m490 net07007 net06997 net09194 vss nmos L=40e-9 W=90e-9
m489 net07067 c14 vss vss nmos L=40e-9 W=90e-9
m488 net07033 c13 vss vss nmos L=40e-9 W=90e-9
m487 net09190 net07068 vss vss nmos L=40e-9 W=90e-9
m486 net09192 net07034 vss vss nmos L=40e-9 W=90e-9
m485 net09194 net06998 vss vss nmos L=40e-9 W=90e-9
m471 net06973 net06966 net09196 vss nmos L=40e-9 W=90e-9
m470 net06942 net06935 net09198 vss nmos L=40e-9 W=90e-9
m469 net06997 c12 vss vss nmos L=40e-9 W=90e-9
m468 net06966 c11 vss vss nmos L=40e-9 W=90e-9
m467 net06935 c10 vss vss nmos L=40e-9 W=90e-9
m466 net09196 net06967 vss vss nmos L=40e-9 W=90e-9
m465 net09198 net06936 vss vss nmos L=40e-9 W=90e-9
m449 net06911 net06904 net09200 vss nmos L=40e-9 W=90e-9
m448 net06880 net06873 net09202 vss nmos L=40e-9 W=90e-9
m447 net06849 net06842 net09204 vss nmos L=40e-9 W=90e-9
m446 net06904 c9 vss vss nmos L=40e-9 W=90e-9
m445 net06873 net08787 vss vss nmos L=40e-9 W=90e-9
m444 net06842 c8 vss vss nmos L=40e-9 W=90e-9
m443 net09200 net06905 vss vss nmos L=40e-9 W=90e-9
m442 net09202 net06874 vss vss nmos L=40e-9 W=90e-9
m441 net09204 net0988 vss vss nmos L=40e-9 W=90e-9
m436 net07105 net07076 net09189 vss nmos L=40e-9 W=90e-9
m435 net07068 net07041 net09191 vss nmos L=40e-9 W=90e-9
m434 net07034 net07007 net09193 vss nmos L=40e-9 W=90e-9
m433 net09189 net07079 vss vss nmos L=40e-9 W=90e-9
m432 net09191 net07044 vss vss nmos L=40e-9 W=90e-9
m431 net09193 net07010 vss vss nmos L=40e-9 W=90e-9
m424 net07079 c14 net09205 vss nmos L=40e-9 W=90e-9
m423 net07044 c13 net09206 vss nmos L=40e-9 W=90e-9
m422 net07010 c12 net09207 vss nmos L=40e-9 W=90e-9
m421 net09205 net07051 vss vss nmos L=40e-9 W=90e-9
m420 net09206 net07017 vss vss nmos L=40e-9 W=90e-9
m419 net09207 net06981 vss vss nmos L=40e-9 W=90e-9
m418 net06998 net06973 net09195 vss nmos L=40e-9 W=90e-9
m417 net06967 net06942 net09197 vss nmos L=40e-9 W=90e-9
m416 net06936 net06911 net09199 vss nmos L=40e-9 W=90e-9
m415 net09195 net06975 vss vss nmos L=40e-9 W=90e-9
m414 net09197 net06944 vss vss nmos L=40e-9 W=90e-9
m413 net09199 net06913 vss vss nmos L=40e-9 W=90e-9
m408 net06975 c11 net09208 vss nmos L=40e-9 W=90e-9
m407 net06944 c10 net09209 vss nmos L=40e-9 W=90e-9
m406 net09208 net06950 vss vss nmos L=40e-9 W=90e-9
m405 net09209 net06919 vss vss nmos L=40e-9 W=90e-9
m404 net06905 net06880 net09201 vss nmos L=40e-9 W=90e-9
m403 net06874 net06849 net09203 vss nmos L=40e-9 W=90e-9
m402 net09201 net06882 vss vss nmos L=40e-9 W=90e-9
m401 net09203 net06851 vss vss nmos L=40e-9 W=90e-9
m394 net06913 c9 net09210 vss nmos L=40e-9 W=90e-9
m393 net06882 net08787 net09211 vss nmos L=40e-9 W=90e-9
m392 net06851 c8 net09212 vss nmos L=40e-9 W=90e-9
m391 net09210 net06888 vss vss nmos L=40e-9 W=90e-9
m390 net09211 net06857 vss vss nmos L=40e-9 W=90e-9
m389 net09212 net0955 vss vss nmos L=40e-9 W=90e-9
m380 net07071 net07064 net09214 vss nmos L=40e-9 W=90e-9
m379 net07036 net07030 net09216 vss nmos L=40e-9 W=90e-9
m378 net07001 net06994 net09218 vss nmos L=40e-9 W=90e-9
m377 net07064 c14 vss vss nmos L=40e-9 W=90e-9
m376 net07030 c13 vss vss nmos L=40e-9 W=90e-9
m375 net09214 net07051 vss vss nmos L=40e-9 W=90e-9
m374 net09216 net07017 vss vss nmos L=40e-9 W=90e-9
m373 net09218 net06981 vss vss nmos L=40e-9 W=90e-9
m366 net07089 net07071 net09213 vss nmos L=40e-9 W=90e-9
m365 net07051 net07036 net09215 vss nmos L=40e-9 W=90e-9
m364 net07017 net07001 net09217 vss nmos L=40e-9 W=90e-9
m363 net09213 net07074 vss vss nmos L=40e-9 W=90e-9
m362 net09215 net07039 vss vss nmos L=40e-9 W=90e-9
m361 net09217 net07004 vss vss nmos L=40e-9 W=90e-9
m354 net07074 c14 net09229 vss nmos L=40e-9 W=90e-9
m353 net07039 c13 net09230 vss nmos L=40e-9 W=90e-9
m352 net07004 c12 net09231 vss nmos L=40e-9 W=90e-9
m351 net09229 net07068 vss vss nmos L=40e-9 W=90e-9
m350 net09230 net07034 vss vss nmos L=40e-9 W=90e-9
m349 net09231 net06998 vss vss nmos L=40e-9 W=90e-9
m341 net06969 net06963 net09220 vss nmos L=40e-9 W=90e-9
m340 net06938 net06932 net09222 vss nmos L=40e-9 W=90e-9
m339 net06994 c12 vss vss nmos L=40e-9 W=90e-9
m338 net06963 c11 vss vss nmos L=40e-9 W=90e-9
m337 net06932 c10 vss vss nmos L=40e-9 W=90e-9
m336 net09220 net06950 vss vss nmos L=40e-9 W=90e-9
m335 net09222 net06919 vss vss nmos L=40e-9 W=90e-9
m328 net06981 net06969 net09219 vss nmos L=40e-9 W=90e-9
m327 net06950 net06938 net09221 vss nmos L=40e-9 W=90e-9
m326 net06919 net06907 net09223 vss nmos L=40e-9 W=90e-9
m325 net09219 net06971 vss vss nmos L=40e-9 W=90e-9
m324 net09221 net06940 vss vss nmos L=40e-9 W=90e-9
m323 net09223 net06909 vss vss nmos L=40e-9 W=90e-9
m318 net06971 c11 net09232 vss nmos L=40e-9 W=90e-9
m317 net06940 c10 net09233 vss nmos L=40e-9 W=90e-9
m316 net09232 net06967 vss vss nmos L=40e-9 W=90e-9
m315 net09233 net06936 vss vss nmos L=40e-9 W=90e-9
m305 net06907 net06901 net09224 vss nmos L=40e-9 W=90e-9
m304 net06876 net06870 net09226 vss nmos L=40e-9 W=90e-9
m303 net06845 net06839 net09228 vss nmos L=40e-9 W=90e-9
m302 net06901 c9 vss vss nmos L=40e-9 W=90e-9
m301 net06870 net08787 vss vss nmos L=40e-9 W=90e-9
m300 net06839 c8 vss vss nmos L=40e-9 W=90e-9
m299 net09224 net06888 vss vss nmos L=40e-9 W=90e-9
m298 net09226 net06857 vss vss nmos L=40e-9 W=90e-9
m297 net09228 net0955 vss vss nmos L=40e-9 W=90e-9
m292 net06888 net06876 net09225 vss nmos L=40e-9 W=90e-9
m291 net06857 net06845 net09227 vss nmos L=40e-9 W=90e-9
m290 net09225 net06878 vss vss nmos L=40e-9 W=90e-9
m289 net09227 net06847 vss vss nmos L=40e-9 W=90e-9
m282 net06909 c9 net09234 vss nmos L=40e-9 W=90e-9
m281 net06878 net08787 net09235 vss nmos L=40e-9 W=90e-9
m280 net06847 c8 net09236 vss nmos L=40e-9 W=90e-9
m279 net09234 net06905 vss vss nmos L=40e-9 W=90e-9
m278 net09235 net06874 vss vss nmos L=40e-9 W=90e-9
m277 net09236 net0988 vss vss nmos L=40e-9 W=90e-9
m241 net0947 net0940 net01050 vss nmos L=40e-9 W=90e-9
m240 net0916 net0909 net01051 vss nmos L=40e-9 W=90e-9
m238 net0940 c7 vss vss nmos L=40e-9 W=90e-9
m237 net0909 c6 vss vss nmos L=40e-9 W=90e-9
m235 net01050 net0941 vss vss nmos L=40e-9 W=90e-9
m234 net01051 net0910 vss vss nmos L=40e-9 W=90e-9
m227 net0988 net0947 net01054 vss nmos L=40e-9 W=90e-9
m226 net0941 net0916 net01056 vss nmos L=40e-9 W=90e-9
m224 net01054 net0949 vss vss nmos L=40e-9 W=90e-9
m223 net01056 net0918 vss vss nmos L=40e-9 W=90e-9
m215 net0949 c7 net01055 vss nmos L=40e-9 W=90e-9
m214 net0918 c6 net01057 vss nmos L=40e-9 W=90e-9
m212 net01055 net0924 vss vss nmos L=40e-9 W=90e-9
m211 net01057 net0893 vss vss nmos L=40e-9 W=90e-9
m200 net0943 net0937 net01063 vss nmos L=40e-9 W=90e-9
m199 net0912 net0906 net01066 vss nmos L=40e-9 W=90e-9
m197 net0937 c7 vss vss nmos L=40e-9 W=90e-9
m196 net0906 c6 vss vss nmos L=40e-9 W=90e-9
m194 net01063 net0924 vss vss nmos L=40e-9 W=90e-9
m193 net01066 net0893 vss vss nmos L=40e-9 W=90e-9
m185 net0955 net0943 net01061 vss nmos L=40e-9 W=90e-9
m184 net0924 net0912 net01064 vss nmos L=40e-9 W=90e-9
m182 net01061 net0945 vss vss nmos L=40e-9 W=90e-9
m181 net01064 net0914 vss vss nmos L=40e-9 W=90e-9
m173 net0945 c7 net01062 vss nmos L=40e-9 W=90e-9
m172 net0914 c6 net01065 vss nmos L=40e-9 W=90e-9
m170 net01062 net0941 vss vss nmos L=40e-9 W=90e-9
m169 net01065 net0910 vss vss nmos L=40e-9 W=90e-9
m161 net0885 net0878 net01069 vss nmos L=40e-9 W=90e-9
m160 net0854 net0847 net01072 vss nmos L=40e-9 W=90e-9
m159 net0878 c5 vss vss nmos L=40e-9 W=90e-9
m158 net0847 c4 vss vss nmos L=40e-9 W=90e-9
m157 net01069 net0879 vss vss nmos L=40e-9 W=90e-9
m156 net01072 net0848 vss vss nmos L=40e-9 W=90e-9
m152 net0910 net0885 net01067 vss nmos L=40e-9 W=90e-9
m151 net0879 net0854 net01070 vss nmos L=40e-9 W=90e-9
m150 net01067 net0887 vss vss nmos L=40e-9 W=90e-9
m149 net01070 net0856 vss vss nmos L=40e-9 W=90e-9
m144 net0887 c5 net01068 vss nmos L=40e-9 W=90e-9
m143 net0856 c4 net01071 vss nmos L=40e-9 W=90e-9
m142 net01068 net0862 vss vss nmos L=40e-9 W=90e-9
m141 net01071 net0831 vss vss nmos L=40e-9 W=90e-9
m134 net0881 net0875 net01075 vss nmos L=40e-9 W=90e-9
m133 net0850 net0844 net01078 vss nmos L=40e-9 W=90e-9
m132 net0875 c5 vss vss nmos L=40e-9 W=90e-9
m131 net0844 c4 vss vss nmos L=40e-9 W=90e-9
m130 net01075 net0862 vss vss nmos L=40e-9 W=90e-9
m129 net01078 net0831 vss vss nmos L=40e-9 W=90e-9
m124 net0893 net0881 net01073 vss nmos L=40e-9 W=90e-9
m123 net0862 net0850 net01076 vss nmos L=40e-9 W=90e-9
m122 net01073 net0883 vss vss nmos L=40e-9 W=90e-9
m121 net01076 net0852 vss vss nmos L=40e-9 W=90e-9
m116 net0883 c5 net01074 vss nmos L=40e-9 W=90e-9
m115 net0852 c4 net01077 vss nmos L=40e-9 W=90e-9
m114 net01074 net0879 vss vss nmos L=40e-9 W=90e-9
m113 net01077 net0848 vss vss nmos L=40e-9 W=90e-9
m108 net0823 net0816 net01081 vss nmos L=40e-9 W=90e-9
m107 net0816 c3 vss vss nmos L=40e-9 W=90e-9
m106 net01081 net0200 vss vss nmos L=40e-9 W=90e-9
m103 net0848 net0823 net01079 vss nmos L=40e-9 W=90e-9
m102 net01079 net0825 vss vss nmos L=40e-9 W=90e-9
m99 net0825 c3 net01080 vss nmos L=40e-9 W=90e-9
m98 net01080 net0198 vss vss nmos L=40e-9 W=90e-9
m94 net0819 net0813 net01084 vss nmos L=40e-9 W=90e-9
m93 net0813 c3 vss vss nmos L=40e-9 W=90e-9
m92 net01084 net0198 vss vss nmos L=40e-9 W=90e-9
m89 net0831 net0819 net01082 vss nmos L=40e-9 W=90e-9
m88 net01082 net0821 vss vss nmos L=40e-9 W=90e-9
m85 net0821 c3 net01083 vss nmos L=40e-9 W=90e-9
m84 net01083 net0200 vss vss nmos L=40e-9 W=90e-9
m80 net0190 net0183 net0227 vss nmos L=40e-9 W=90e-9
m79 net0183 c2 vss vss nmos L=40e-9 W=90e-9
m78 net0227 net55 vss vss nmos L=40e-9 W=90e-9
m75 net0200 net0190 net0226 vss nmos L=40e-9 W=90e-9
m74 net0226 net0192 vss vss nmos L=40e-9 W=90e-9
m71 net0192 c2 net0228 vss nmos L=40e-9 W=90e-9
m70 net0228 net51 vss vss nmos L=40e-9 W=90e-9
m66 net0186 net0180 net0231 vss nmos L=40e-9 W=90e-9
m65 net0180 c2 vss vss nmos L=40e-9 W=90e-9
m64 net0231 net51 vss vss nmos L=40e-9 W=90e-9
m61 net0198 net0186 net0229 vss nmos L=40e-9 W=90e-9
m60 net0229 net0188 vss vss nmos L=40e-9 W=90e-9
m57 net0188 c2 net0230 vss nmos L=40e-9 W=90e-9
m56 net0230 net55 vss vss nmos L=40e-9 W=90e-9
m27 net168 net32 vss vss nmos L=40e-9 W=90e-9
m26 net51 net28 net168 vss nmos L=40e-9 W=90e-9
m23 net169 start1 vss vss nmos L=40e-9 W=90e-9
m22 net32 c1 net169 vss nmos L=40e-9 W=90e-9
m19 net19 c1 vss vss nmos L=40e-9 W=90e-9
m17 net170 start2 vss vss nmos L=40e-9 W=90e-9
m16 net28 net19 net170 vss nmos L=40e-9 W=90e-9
m13 net171 net39 vss vss nmos L=40e-9 W=90e-9
m12 net55 net36 net171 vss nmos L=40e-9 W=90e-9
m9 net172 start2 vss vss nmos L=40e-9 W=90e-9
m8 net39 c1 net172 vss nmos L=40e-9 W=90e-9
m5 net22 c1 vss vss nmos L=40e-9 W=90e-9
m0 net173 start1 vss vss nmos L=40e-9 W=90e-9
m2 net36 net22 net173 vss nmos L=40e-9 W=90e-9
xi11 net03559 net03557 out vdd vss Arbiter
xi10 net04550 net04530 net05098 vdd vss Arbiter
xi8 net08576 net08559 net08884 vdd vss Arbiter
xi7 net08295 net08278 net08868 vdd vss Arbiter
xi6 net08014 net07997 net08852 vdd vss Arbiter
xi5 net07733 net07716 net08836 vdd vss Arbiter
xi4 net07449 net07432 net08819 vdd vss Arbiter
xi3 net07167 net07150 net08803 vdd vss Arbiter
xi2 net06874 net06857 net08787 vdd vss Arbiter

