** Generated for: hspiceD
** Generated on: Jun 14 12:58:44 2013
** Design library name: FFPUF_SCA
** Design cell name: 128stagesMux2Arb
** Design view name: schematic
.GLOBAL vss! vdd!

.include '/home/akommini/658proj/NMOS32LP.inc'
.include '/home/akommini/658proj/PMOS32LP.inc'
vsupply vdd! 0 1.0
vss vss! 0 0
.vec '68stage2FFPUF1.vec'
vclock clk 0 PWL (0 0 3.49n 0 3.5n 1.1 3.9n 1.1)

.TEMP 25
.OPTION
+ POST=2
+ PROBE

** Library name: NangateOpenCellLibrary
** Cell name: NAND2_X1
** View name: schematic
.subckt NAND2_X1 a1 a2 zn
m_i_3 zn a2 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9
m_i_2 vdd! a1 zn vdd! PMOS_VTL L=50e-9 W=630e-9
m_i_0 zn a1 net_0 vss! NMOS_VTL L=50e-9 W=415e-9
m_i_1 net_0 a2 vss! vss! NMOS_VTL L=50e-9 W=415e-9
.ends NAND2_X1
** End of subcircuit definition.

** Library name: NangateOpenCellLibrary
** Cell name: INV_X1
** View name: schematic
.subckt INV_X1 a zn
m_i_0 zn a vss! vss! NMOS_VTL L=50e-9 W=415e-9
m_i_1 zn a vdd! vdd! PMOS_VTL L=50e-9 W=630e-9
.ends INV_X1
** End of subcircuit definition.

** Library name: FFPUF_SCA
** Cell name: Arbiter
** View name: schematic
.subckt Arbiter a b y_a y_b
xi1 net6 b net5 NAND2_X1
xi0 net5 a net6 NAND2_X1
xi5 net5 y_b INV_X1
xi4 net6 y_a INV_X1
.ends Arbiter
** End of subcircuit definition.

** Library name: NangateOpenCellLibrary
** Cell name: DFF_X1
** View name: schematic
.subckt DFF_X1 ck d q qn
m_mn3 z2 d vss! vss! NMOS_VTL L=50e-9 W=275e-9
m_mn4 z2 cni z3 vss! NMOS_VTL L=50e-9 W=275e-9
m_mn6 vss! z4 z6 vss! NMOS_VTL L=50e-9 W=90e-9
m_mn7 z3 ci z6 vss! NMOS_VTL L=50e-9 W=90e-9
m_mn1 vss! ck cni vss! NMOS_VTL L=50e-9 W=210e-9
m_mn8 z12 z3 vss! vss! NMOS_VTL L=50e-9 W=210e-9
m_mn9 z9 ci z12 vss! NMOS_VTL L=50e-9 W=210e-9
m_mn12 z9 cni z8 vss! NMOS_VTL L=50e-9 W=90e-9
m_mn11 z8 z10 vss! vss! NMOS_VTL L=50e-9 W=90e-9
m_mn14 qn z9 vss! vss! NMOS_VTL L=50e-9 W=415e-9
m_mn13 vss! z10 q vss! NMOS_VTL L=50e-9 W=415e-9
m_mn5 z4 z3 vss! vss! NMOS_VTL L=50e-9 W=210e-9
m_mn2 ci cni vss! vss! NMOS_VTL L=50e-9 W=210e-9
m_mn10 vss! z9 z10 vss! NMOS_VTL L=50e-9 W=210e-9
m_mp4 z3 ci z5 vdd! PMOS_VTL L=50e-9 W=420e-9
m_mp3 z5 d vdd! vdd! PMOS_VTL L=50e-9 W=420e-9
m_mp7 z1 cni z3 vdd! PMOS_VTL L=50e-9 W=90e-9
m_mp6 vdd! z4 z1 vdd! PMOS_VTL L=50e-9 W=90e-9
m_mp1 vdd! ck cni vdd! PMOS_VTL L=50e-9 W=315e-9
m_mp8 z7 z3 vdd! vdd! PMOS_VTL L=50e-9 W=315e-9
m_mp9 z9 cni z7 vdd! PMOS_VTL L=50e-9 W=315e-9
m_mp12 z9 ci z11 vdd! PMOS_VTL L=50e-9 W=90e-9
m_mp11 z11 z10 vdd! vdd! PMOS_VTL L=50e-9 W=90e-9
m_mp14 qn z9 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9
m_mp13 vdd! z10 q vdd! PMOS_VTL L=50e-9 W=630e-9
m_mp5 z4 z3 vdd! vdd! PMOS_VTL L=50e-9 W=315e-9
m_mp2 ci cni vdd! vdd! PMOS_VTL L=50e-9 W=315e-9
m_mp10 vdd! z9 z10 vdd! PMOS_VTL L=50e-9 W=315e-9
.ends DFF_X1
** End of subcircuit definition.

** Library name: FFPUF_SCA
** Cell name: 128stagesMux2Arb
** View name: schematic
m3154 s128a net028885 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.064818
m3152 net028885 net028897 net022149 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.000386
m3151 net022149 s127a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.044414
m3148 vss! chal128 net028897 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.060083
m3147 s127a net028921 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.033654
m3145 net028921 net028933 net022165 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.104280
m3144 net022165 s126a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.044057
m3143 vss! chal127 net028933 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.041577
m3140 s126a net028965 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.044009
m3138 net028965 net028945 net022181 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.024938
m3137 net022181 s125a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.091356
m3134 vss! chal126 net028945 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.025597
m3133 net022197 s124a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.054045
m3132 net21589 net029005 net022197 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.087873
m3131 s125a net21589 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.008983
m3129 vss! chal125 net029005 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.066404
m3125 net022213 s123a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.008715
m3124 net029037 net029033 net022213 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.146996
m3123 s124a net029037 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.018220
m3122 vss! chal124 net029033 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.038184
m3118 s123a net029065 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.007030
m3115 vss! chal123 net029077 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.051303
m3114 net029065 net029077 net022233 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.106691
m3113 net022233 s122a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.024485
m3110 net029101 net029113 net022241 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.016300
m3109 net022241 s121a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.045780
m3108 s122a net029101 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.059147
m3106 vss! chal122 net029113 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.056358
m3105 net022261 s120a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.034353
m3104 net029145 net029141 net022261 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.070400
m3103 s121a net029145 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.188395
m3101 vss! chal121 net029141 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.026007
m3098 s120a net029173 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.045719
m3096 net029173 net029185 net022277 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.029703
m3095 net022277 s119a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.086067
m3092 vss! chal120 net029185 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.047432
m3091 s119a net029209 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.064165
m3089 net029209 net029221 net022293 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.033652
m3088 net022293 s118a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.105500
m3087 vss! chal119 net029221 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.053193
m3084 s118a net029245 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.074189
m3082 net029245 net029257 net022309 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.013866
m3080 net022309 s117a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.018144
m3078 vss! chal118 net029257 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.038845
m3077 net20711 net029293 net022321 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.071500
m3076 s117a net20711 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.013308
m3074 net022321 s116a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.030435
m3073 vss! chal117 net029293 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.103192
m3068 s116a net029317 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.027526
m3067 net029317 net029329 net022341 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.059086
m3066 net022341 s115a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.035198
m3064 vss! chal116 net029329 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.093745
m3063 net022357 s114a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.042207
m3062 net029361 net029357 net022357 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.030767
m3061 s115a net029361 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.110005
m3059 vss! chal115 net029357 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.079208
m3055 s114a net029389 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.024172
m3054 net022377 s113a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.036637
m3053 net029389 net029401 net022377 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.073077
m3052 vss! chal114 net029401 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.088191
m3048 s113a net029425 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.077412
m3045 net029425 net029437 net022389 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.004296
m3044 net022389 s112a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.086149
m3043 vss! chal113 net029437 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.038157
m3041 s112a net029469 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.097998
m3038 vss! chal112 net029465 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.085154
m3037 net022413 s111a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.164066
m3036 net029469 net029465 net022413 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.183402
m3033 net022421 s110a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.023230
m3032 net029497 net029509 net022421 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.023704
m3030 s111a net029497 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.099654
m3029 vss! chal111 net029509 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.036487
m3027 s110a net029533 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.099556
m3024 net022441 s109a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.004151
m3023 net029533 net029545 net022441 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.067241
m3022 vss! chal110 net029545 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.114444
m3018 s109a net19022 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.020319
m3017 net19022 net029581 net022453 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.028673
m3016 net022453 s108a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.092198
m3015 vss! chal109 net029581 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.019411
m3012 s108a net029609 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.050028
m3011 net029609 net029613 net022469 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.015350
m3010 net022469 s107a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.015791
m3008 vss! chal108 net029613 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.050985
m3007 s107a net029641 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.080128
m3005 vss! chal107 net029653 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.026438
m3002 net022493 s106a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.001024
m3001 net029641 net029653 net022493 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.062697
m2999 s106a net029677 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.024657
m2998 net022505 s105a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.010089
m2997 net029677 net029689 net022505 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.018246
m2996 vss! chal106 net029689 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.063821
m2992 s105a net029717 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.161433
m2991 net029717 net029721 net022517 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.059335
m2990 net022517 s104a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.044988
m2987 vss! chal105 net029721 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.000330
m2985 s104a net029749 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.009085
m2982 vss! chal104 net029761 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.040700
m2981 net022541 s103a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.038709
m2980 net029749 net029761 net022541 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.104479
m2977 net022549 s102a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.030038
m2976 net029785 net029797 net022549 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.049131
m2974 s103a net029785 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.027560
m2973 vss! chal103 net029797 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.058138
m2971 s102a net029821 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.087739
m2968 net022569 s101a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.098240
m2967 net029821 net029833 net022569 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.019677
m2966 vss! chal102 net029833 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.136818
m2962 s101a net19841 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.014031
m2961 net19841 net029861 net022581 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.034335
m2960 net022581 s100a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.010067
m2959 vss! chal101 net029861 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.016107
m2957 s100a net029893 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.165583
m2956 net022601 s99a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.054689
m2955 net029893 net029905 net022601 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.011122
m2952 vss! chal100 net029905 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.047160
m2950 s99a net029933 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.049983
m2949 net029933 net029937 net022613 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.017863
m2948 net022613 s98a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.022908
m2945 vss! chal99 net029937 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.051947
m2944 s98a net029965 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.070399
m2943 net029965 net029977 net022629 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.008359
m2942 net022629 s97a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.014031
m2938 vss! chal98 net029977 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.110170
m2937 s97a net030009 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.037704
m2935 net022649 s96a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.002314
m2934 net030009 net030005 net022649 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.093922
m2931 vss! chal97 net030005 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.102964
m2930 s96a net030045 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.041344
m2928 net030045 net030025 net022661 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.049013
m2927 net022661 s95a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.016883
m2926 vss! chal96 net030025 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.060859
m2923 s95a net030073 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.012712
m2921 net030073 net030085 net022677 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.015952
m2920 net022677 s94a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.122130
m2917 vss! chal95 net030085 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.127251
m2916 s94a net030109 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.074314
m2915 net030109 net030121 net022693 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.075879
m2914 net022693 s93a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.081877
m2912 vss! chal94 net030121 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.089304
m2909 s93a net20343 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.065910
m2907 net022713 s92a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.111962
m2906 net20343 net030157 net022713 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.221638
m2903 vss! chal93 net030157 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.022307
m2899 s92a net030181 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.046406
m2898 net022729 s91a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.000555
m2897 net030181 net030193 net022729 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.004831
m2896 vss! chal92 net030193 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.144902
m2894 net022741 s90a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.050089
m2893 net030217 net030229 net022741 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.037052
m2892 s91a net030217 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.002488
m2889 vss! chal91 net030229 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.116403
m2887 s90a net030261 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.034404
m2884 net022761 s89a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.010505
m2883 net030261 net030257 net022761 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.005693
m2882 vss! chal90 net030257 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.117514
m2880 net022773 s88a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.017874
m2879 net030297 net030277 net022773 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.107034
m2878 s89a net030297 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.111491
m2877 vss! chal89 net030277 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.030715
m2873 s88a net030325 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.094056
m2870 net030325 net030337 net022789 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.026624
m2869 net022789 s87a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.041234
m2868 vss! chal88 net030337 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.033253
m2866 s87a net030361 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.012963
m2865 net030361 net030373 net022805 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.080130
m2864 net022805 s86a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.008505
m2861 vss! chal87 net030373 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.038683
m2859 s86a net030397 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.046062
m2856 net022825 s85a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.101308
m2855 net030397 net030409 net022825 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.008194
m2854 vss! chal86 net030409 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.044095
m2852 s85a net030437 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.026272
m2851 net030437 net030441 net022837 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.071042
m2850 net022837 s84a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.132290
m2847 vss! chal85 net030441 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.100363
m2845 s84a net030469 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.019316
m2842 net022857 s83a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.021085
m2841 net030469 net030481 net022857 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.053165
m2840 vss! chal84 net030481 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.026596
m2838 net022869 s82a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.092561
m2837 net030505 net030517 net022869 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.006743
m2836 s83a net030505 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.077073
m2833 vss! chal83 net030517 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.018579
m2831 s82a net030541 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.013017
m2830 vss! chal82 net030553 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.029465
m2827 net022893 s81a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.088769
m2826 net030541 net030553 net022893 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.064002
m2824 s81a net19306 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.030076
m2823 net19306 net030589 net022901 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.094248
m2822 net022901 s80a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.063949
m2820 vss! chal81 net030589 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.023333
m2818 s128b net028869 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.076481
m2816 net022914 s127a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.027087
m2814 net028869 net028893 net022921 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.008570
m2813 net028869 chal128 net022914 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.046184
m2810 net022921 s127b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.043713
m2808 net022930 s127b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.015842
m2806 net028885 chal128 net022930 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.038559
m2803 vss! chal128 net028893 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.093959
m2801 net022942 s126a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.051561
m2800 s127b net028905 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.064368
m2799 net028905 net028929 net022953 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.072453
m2798 net028905 chal127 net022942 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.024039
m2796 net022953 s126b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.021552
m2795 net022962 s126b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.090690
m2794 net028921 chal127 net022962 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.018276
m2786 vss! chal127 net028929 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.028159
m2784 s126b net028949 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.057887
m2782 net022978 s125a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.036205
m2781 net028949 chal126 net022978 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.027994
m2780 net022993 s125b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.059299
m2779 net028949 net028941 net022993 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.003361
m2778 net022994 s125b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.034505
m2777 net028965 chal126 net022994 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.023481
m2775 vss! chal126 net028941 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.046985
m2767 s125b net028977 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.029516
m2765 net023010 s124a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.101019
m2763 net028977 chal125 net023010 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.025500
m2761 net028977 net15878 net17576 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.062880
m2760 net17576 s124b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.067784
m2757 net19531 s124b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.003964
m2755 net21589 chal125 net19531 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.005927
m2752 vss! chal125 net15878 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.061041
m2750 s124b net029021 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.126256
m2748 net023042 s123a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.002362
m2747 net029021 chal124 net023042 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.004840
m2746 net029021 net029013 net023053 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.025591
m2745 net023053 s123b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.061940
m2744 net023058 s123b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.098712
m2743 net029037 chal124 net023058 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.184687
m2738 vss! chal124 net029013 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.038157
m2733 s123b net029049 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.075460
m2729 net029049 chal123 net023078 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.031103
m2728 net023078 s122a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.166553
m2726 net029049 net029073 net023085 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.044868
m2724 net023085 s122b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.091790
m2722 net023090 s122b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.010198
m2720 net029065 chal123 net023090 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.007405
m2718 vss! chal123 net029073 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.047765
m2716 net023102 s121a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.008473
m2715 net029085 net029109 net023109 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.053453
m2714 net029085 chal122 net023102 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.106612
m2713 net023109 s121b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.041069
m2712 net023118 s121b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.095462
m2711 net029101 chal122 net023118 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.050652
m2710 s122b net029085 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.007254
m2701 vss! chal122 net029109 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.129710
m2699 s121b net029125 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.025592
m2697 net023138 s120a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.064569
m2696 net029125 chal121 net023138 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.094526
m2695 net029125 net029121 net023149 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.003654
m2694 net023149 s120b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.016046
m2693 net023154 s120b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.055117
m2692 net029145 chal121 net023154 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.036611
m2688 vss! chal121 net029121 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.004543
m2682 s120b net029157 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.015132
m2680 net023170 s119a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.022419
m2678 net029157 chal120 net023170 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.045037
m2676 net023185 s119b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.170744
m2675 net029157 net029181 net023185 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.011598
m2672 net023186 s119b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.073374
m2670 net029173 chal120 net023186 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.013347
m2667 vss! chal120 net029181 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.040469
m2665 s119b net029193 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.041685
m2663 net023202 s118a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.012092
m2661 net029193 chal119 net023202 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.040878
m2659 net023217 s118b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.080152
m2658 net029193 net029217 net023217 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.032896
m2655 net023218 s118b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.096315
m2653 net029209 chal119 net023218 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.002923
m2650 vss! chal119 net029217 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.004152
m2648 s118b net029229 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.021931
m2646 net023234 s117a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.101387
m2644 net029229 chal118 net023234 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.167310
m2642 net023249 s117b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.117359
m2641 net029229 net029253 net023249 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.088673
m2638 net023250 s117b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.132547
m2636 net029245 chal118 net023250 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.014334
m2633 vss! chal118 net029253 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.094767
m2631 net023262 s116a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.151914
m2630 net029265 chal117 net023262 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.013279
m2629 s117b net029265 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.031887
m2628 net029265 net16859 net18435 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.033404
m2627 net18435 s116b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.017929
m2625 net19505 s116b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.055907
m2624 net20711 chal117 net19505 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.011945
m2616 vss! chal117 net16859 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.142612
m2614 net029301 chal116 net023298 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.023778
m2613 net023298 s115a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.050110
m2612 net029301 net029325 net023305 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.038116
m2611 s116b net029301 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.016472
m2610 net023305 s115b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.032377
m2608 net023314 s115b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.146571
m2607 net029317 chal116 net023314 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.010500
m2599 vss! chal116 net029325 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.128347
m2597 s115b net029345 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.012974
m2595 net023330 s114a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.053549
m2594 net029345 chal115 net023330 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.082571
m2593 net029345 net029337 net023341 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.052708
m2592 net023341 s114b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.033885
m2591 net023346 s114b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.054281
m2590 net029361 chal115 net023346 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.003966
m2585 vss! chal115 net029337 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.002695
m2580 s114b net029377 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.071431
m2578 net023362 s113a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.076110
m2577 net029377 chal114 net023362 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.032958
m2574 net029377 net029397 net023373 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.125810
m2572 net023373 s113b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.160673
m2570 net023378 s113b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.113581
m2568 net029389 chal114 net023378 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.070005
m2565 vss! chal114 net029397 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.031298
m2563 net029409 chal113 net023394 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.054309
m2562 net023394 s112a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.005973
m2561 s113b net029409 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.025857
m2560 net029409 net029433 net023405 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.097035
m2558 net023405 s112b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.059517
m2557 net023410 s112b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.052457
m2556 net029425 chal113 net023410 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.056125
m2548 vss! chal113 net029433 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.030747
m2546 s112b net029453 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.055103
m2544 net023426 s111a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.035523
m2543 net029453 chal112 net023426 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.048602
m2542 net029453 net029445 net023437 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.023823
m2541 net023437 s111b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.013430
m2540 net023442 s111b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.068252
m2539 net029469 chal112 net023442 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.149811
m2533 vss! chal112 net029445 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.102713
m2529 s111b net029485 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.110882
m2521 net023458 s110a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.037094
m2520 net029485 chal111 net023458 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.087279
m2519 net029485 net029505 net023469 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.140756
m2518 net023469 s110b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.084750
m2517 net023474 s110b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.152734
m2516 net029497 chal111 net023474 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.079189
m2514 vss! chal111 net029505 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.094801
m2512 s110b net029517 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.033354
m2509 net023490 s109a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.187651
m2506 net029517 chal110 net023490 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.027357
m2505 net029517 net029541 net023501 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.070280
m2503 net023501 s109b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.010220
m2501 net023506 s109b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.019570
m2499 net029533 chal110 net023506 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.054836
m2497 vss! chal110 net029541 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.011257
m2495 s109b net029553 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.103805
m2492 net023522 s108a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.059505
m2489 net029553 net16774 net17356 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.074846
m2488 net029553 chal109 net023522 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.011784
m2486 net17356 s108b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.106113
m2484 net19023 s108b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.151027
m2482 net19022 chal109 net19023 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.122899
m2480 vss! chal109 net16774 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.024272
m2478 s108b net029589 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.045787
m2476 net029589 chal108 net023558 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.075703
m2475 net023558 s107a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.007237
m2474 net029589 net029597 net023565 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.033031
m2473 net023565 s107b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.003578
m2472 net023570 s107b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.053795
m2471 net029609 chal108 net023570 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.065484
m2465 vss! chal108 net029597 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.010690
m2461 s107b net029629 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.119025
m2453 net023586 s106a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.026828
m2452 net029629 chal107 net023586 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.069220
m2451 net029629 net029649 net023597 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.122199
m2450 net023597 s106b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.027360
m2449 net023602 s106b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.094640
m2448 net029641 chal107 net023602 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.015330
m2446 vss! chal107 net029649 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.031520
m2444 net023614 s105a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.019497
m2443 net029665 chal106 net023614 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.112272
m2442 s106b net029665 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.063775
m2441 net029665 net029685 net023629 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.013511
m2439 net023629 s105b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.005018
m2438 net023634 s105b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.013392
m2437 net029677 chal106 net023634 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.044886
m2429 vss! chal106 net029685 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.092999
m2427 s105b net029697 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.013612
m2425 net029697 chal105 net023654 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.054313
m2424 net023654 s104a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.053105
m2423 net029697 net029705 net023661 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.005292
m2422 net023661 s104b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.065030
m2421 net023666 s104b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.029720
m2420 net029717 chal105 net023666 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.061010
m2414 vss! chal105 net029705 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.015857
m2410 s104b net029737 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.039433
m2406 net023682 s103a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.057206
m2405 net029737 chal104 net023682 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.012414
m2403 net029737 net029757 net023693 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.007233
m2401 net023693 s103b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.063349
m2399 net023698 s103b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.055604
m2397 net029749 chal104 net023698 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.037739
m2395 vss! chal104 net029757 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.036516
m2393 s103b net029769 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.021798
m2390 net023714 s102a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.057829
m2387 net029769 chal103 net023714 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.024496
m2386 net029769 net029793 net023725 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.008085
m2384 net023725 s102b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.086438
m2382 net023730 s102b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.037794
m2380 net029785 chal103 net023730 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.143007
m2378 vss! chal103 net029793 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.090222
m2376 net023742 s101a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.020359
m2375 s102b net029805 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.015105
m2374 net029805 chal102 net023742 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.192594
m2373 net029805 net029829 net023757 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.099055
m2371 net023757 s101b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.017071
m2370 net023762 s101b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.002818
m2369 net029821 chal102 net023762 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.096168
m2361 vss! chal102 net029829 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.075543
m2359 s101b net029841 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.052075
m2357 net023778 s100a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.108000
m2356 net029841 net16703 net17250 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.048127
m2355 net029841 chal101 net023778 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.248512
m2354 net17250 s100b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.067694
m2353 net19424 s100b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.021825
m2352 net19841 chal101 net19424 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.057055
m2346 vss! chal101 net16703 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.019836
m2342 net023806 s99a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.004637
m2341 net029881 chal100 net023806 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.038325
m2340 net029881 net029901 net023817 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.004764
m2339 net023817 s99b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.035908
m2338 net023822 s99b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.080017
m2337 net029893 chal100 net023822 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.062576
m2336 s100b net029881 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.040024
m2327 vss! chal100 net029901 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.050445
m2325 s99b net029913 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.059353
m2323 net029913 chal99 net023846 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.110084
m2322 net023846 s98a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.073900
m2321 net029913 net029921 net023853 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.093871
m2320 net023853 s98b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.017449
m2319 net023858 s98b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.056119
m2318 net029933 chal99 net023858 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.047582
m2313 vss! chal99 net029921 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.120847
m2308 net029949 chal98 net023874 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.035424
m2307 net023874 s97a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.065045
m2306 net029949 net029973 net023881 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.108045
m2305 s98b net029949 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.039974
m2304 net023881 s97b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.010775
m2302 net023890 s97b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.038733
m2301 net029965 chal98 net023890 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.089375
m2293 vss! chal98 net029973 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.044759
m2291 net023902 s96a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.105415
m2290 net029993 chal97 net023902 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.066038
m2289 s97b net029993 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.002858
m2288 net029993 net029985 net023917 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.021487
m2287 net023917 s96b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.074678
m2285 net023922 s96b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.022620
m2284 net030009 chal97 net023922 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.065511
m2279 vss! chal97 net029985 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.099163
m2274 s96b net030029 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.025385
m2272 net030029 chal96 net023942 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.133957
m2271 net023942 s95a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.022395
m2270 net030029 net030021 net023949 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.119041
m2269 net023949 s95b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.055364
m2268 net023954 s95b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.097102
m2267 net030045 chal96 net023954 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.012794
m2265 vss! chal96 net030021 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.063588
m2257 s95b net030057 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.085885
m2255 net030057 chal95 net023974 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.035749
m2254 net023974 s94a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.057293
m2251 net030057 net030081 net023981 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.088324
m2249 net023981 s94b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.102735
m2247 net023986 s94b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.019305
m2245 net030073 chal95 net023986 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.023222
m2242 vss! chal95 net030081 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.055194
m2240 s94b net030093 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.003969
m2238 net030093 chal94 net024006 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.014678
m2237 net024006 s93a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.120503
m2234 net030093 net030117 net024013 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.054282
m2232 net024013 s93b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.007310
m2230 net024018 s93b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.029970
m2228 net030109 chal94 net024018 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.089253
m2225 vss! chal94 net030117 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.128200
m2223 net024030 s92a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.012684
m2222 net030133 chal93 net024030 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.008020
m2221 net030133 net16587 net16590 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.050565
m2220 net16590 s92b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.007840
m2219 net19383 s92b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.116289
m2218 net20343 chal93 net19383 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.073527
m2217 s93b net030133 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.024562
m2208 vss! chal93 net16587 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.099336
m2206 s92b net030169 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.050956
m2202 net024066 s91a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.084424
m2201 net030169 chal92 net024066 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.060074
m2199 net030169 net030189 net024077 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.099607
m2197 net024077 s91b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.057639
m2195 net024082 s91b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.052918
m2193 net030181 chal92 net024082 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.071158
m2191 vss! chal92 net030189 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.046137
m2189 net024094 s90a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.007422
m2188 net030205 chal91 net024094 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.128406
m2187 s91b net030205 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.158001
m2186 net030205 net030225 net024109 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.031021
m2184 net024109 s90b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.002101
m2183 net024114 s90b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.072736
m2182 net030217 chal91 net024114 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.042526
m2174 vss! chal91 net030225 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.016312
m2172 s90b net030245 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.014663
m2170 net024130 s89a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.054882
m2169 net030245 chal90 net024130 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.159039
m2168 net030245 net030237 net024141 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.010966
m2167 net024141 s89b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.083851
m2166 net024146 s89b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.015956
m2165 net030261 chal90 net024146 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.172781
m2159 vss! chal90 net030237 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.002372
m2155 s89b net030285 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.105667
m2153 net024162 s88a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.077750
m2152 net030285 chal89 net024162 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.089290
m2151 net030285 net030273 net024173 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.117153
m2150 net024173 s88b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.019595
m2149 net024178 s88b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.020353
m2148 net030297 chal89 net024178 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.043407
m2146 vss! chal89 net030273 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.008698
m2138 s88b net030309 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.075756
m2134 net030309 chal88 net024198 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.085237
m2133 net024198 s87a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.050551
m2131 net030309 net030333 net024205 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.071342
m2129 net024205 s87b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.040536
m2127 net024210 s87b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.066537
m2125 net030325 chal88 net024210 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.086944
m2123 vss! chal88 net030333 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.018894
m2121 s87b net030345 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.019843
m2118 net024226 s86a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.058729
m2115 net030345 net030369 net024233 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.019377
m2114 net030345 chal87 net024226 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.022611
m2112 net024233 s86b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.065523
m2110 net024242 s86b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.083242
m2108 net030361 chal87 net024242 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.135445
m2106 vss! chal87 net030369 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.061096
m2104 net024254 s85a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.070850
m2103 net030381 chal86 net024254 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.003272
m2102 net030381 net030405 net024265 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.005818
m2101 net024265 s85b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.006385
m2100 net024270 s85b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.044674
m2099 net030397 chal86 net024270 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.015845
m2098 s86b net030381 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.021484
m2089 vss! chal86 net030405 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.094470
m2087 s85b net030417 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.080933
m2085 net024290 s84a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.014414
m2084 net030417 net030421 net024297 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.074648
m2083 net030417 chal85 net024290 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.029475
m2082 net024297 s84b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.076175
m2081 net024306 s84b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.055521
m2080 net030437 chal85 net024306 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.189129
m2074 vss! chal85 net030421 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.034481
m2069 s84b net030453 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.109742
m2067 net024322 s83a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.034892
m2065 net030453 chal84 net024322 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.055413
m2062 net030453 net030477 net024333 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.006507
m2061 net024333 s83b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.026615
m2059 net024338 s83b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.048714
m2057 net030469 chal84 net024338 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.162194
m2055 vss! chal84 net030477 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.018788
m2052 s83b net030489 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.100591
m2050 net024354 s82a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.037751
m2048 net030489 chal83 net024354 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.030105
m2045 net030489 net030513 net024365 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.045551
m2044 net024365 s82b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.063144
m2042 net024370 s82b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.065959
m2040 net030505 chal83 net024370 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.117829
m2038 vss! chal83 net030513 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.169452
m2035 s82b net030525 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.011124
m2033 net024386 s81a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.023022
m2031 net030525 chal82 net024386 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.089278
m2028 net030525 net030549 net024397 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.008377
m2027 net024397 s81b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.066810
m2025 net024402 s81b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.016839
m2023 net030541 chal82 net024402 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.047565
m2021 vss! chal82 net030549 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.067814
m2019 net024414 s80a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.005348
m2018 net030561 chal81 net024414 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.041845
m2016 net16981 s80b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.016589
m2015 net030561 net15612 net16981 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.160766
m2014 s81b net030561 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.098291
m2013 net19304 s80b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.002392
m2012 net19306 chal81 net19304 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.022463
m2004 vss! chal81 net15612 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.026557
m1906 net015276 s79a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.125488
m1904 net019119 chal80 net015276 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.063862
m1900 s80b net019119 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.045984
m1899 net019119 net019159 net015291 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.100364
m1898 net015291 s79b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.059360
m1895 net015296 s79b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.069448
m1894 net019139 chal80 net015296 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.050068
m1892 s80a net019139 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.032575
m1891 net019139 net019163 net015311 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.106571
m1888 net015311 s79a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.108937
m1886 vss! chal80 net019159 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.007197
m1884 vss! chal80 net019163 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.016386
m1883 net015324 s78a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.056548
m1882 net019179 chal79 net015324 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.056435
m1880 s79b net019179 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.017442
m1879 net019179 net019175 net015339 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.077163
m1878 net015339 s78b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.025712
m1877 net019199 chal79 net015348 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.077000
m1876 net015348 s78b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.018443
m1875 net019199 net019195 net015355 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.013376
m1874 s79a net019199 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.122412
m1872 net015355 s78a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.054824
m1866 vss! chal79 net019175 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.044316
m1861 vss! chal79 net019195 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.141567
m1858 s78b net019227 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.028934
m1857 s78a net019247 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.044425
m1853 net015380 s77a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.022369
m1851 net019227 chal78 net015380 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.024377
m1848 vss! chal78 net019223 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.000249
m1847 net019227 net019223 net015395 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.043245
m1846 net015395 s77b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.162994
m1842 net019247 chal78 net015404 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.062050
m1841 net015404 s77b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.017086
m1839 vss! chal78 net019243 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.138119
m1838 net019247 net019243 net015415 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.017434
m1836 net015415 s77a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.018268
m1834 s77b net019279 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.055404
m1833 s77a net019295 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.070653
m1830 vss! chal77 net019271 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.027361
m1828 vss! chal77 net019275 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.041083
m1826 net015436 s76a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.034033
m1824 net019279 chal77 net015436 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.047870
m1821 net019279 net019271 net015447 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.032720
m1820 net015447 s76b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.077741
m1817 net019295 chal77 net015456 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.036578
m1816 net015456 s76b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.050879
m1814 net019295 net019275 net015463 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.157874
m1812 net015463 s76a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.124038
m1809 net015468 s75a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.001861
m1807 net019311 chal76 net015468 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.022995
m1804 net019311 net019315 net015479 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.066418
m1803 s76b net019311 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.037551
m1802 vss! chal76 net019315 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.088132
m1800 net015479 s75b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.047862
m1796 net015492 s75b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.109438
m1795 net019339 chal76 net015492 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.051139
m1793 s76a net019339 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.059767
m1792 net019339 net019343 net015507 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.023713
m1791 vss! chal76 net019343 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.046990
m1788 net015507 s75a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.058913
m1786 net015516 s74a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.133694
m1784 net019359 chal75 net015516 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.023308
m1781 net019359 net019399 net015527 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.010670
m1780 s75b net019359 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.020045
m1778 net015527 s74b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.121256
m1775 net015536 s74b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.079914
m1774 net019383 chal75 net015536 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.032891
m1772 s75a net019383 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.024597
m1771 net019383 net019403 net015551 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.081271
m1768 net015551 s74a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.078796
m1766 vss! chal75 net019399 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.004672
m1764 vss! chal75 net019403 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.009918
m1762 net015564 s73a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.007650
m1760 net019407 chal74 net015564 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.038498
m1758 net019407 net019447 net015575 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.128190
m1756 net015575 s73b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.009161
m1753 net019423 chal74 net015584 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.109548
m1752 net015584 s73b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.011527
m1750 net019423 net019451 net015591 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.014514
m1748 net015591 s73a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.013857
m1747 s74b net019407 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.097039
m1745 s74a net019423 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.025662
m1742 vss! chal74 net019447 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.084733
m1740 vss! chal74 net019451 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.017617
m1739 net015612 s72a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.042224
m1738 net019463 chal73 net015612 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.111888
m1737 net019463 net019467 net015623 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.143556
m1736 s73b net019463 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.058048
m1734 net015623 s72b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.011351
m1733 net015632 s72b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.005272
m1732 net019487 chal73 net015632 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.039368
m1731 s73a net019487 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.016391
m1730 net019487 net019491 net015647 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.018103
m1728 net015647 s72a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.043313
m1723 vss! chal73 net019467 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.037702
m1716 vss! chal73 net019491 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.043140
m1715 s72b net019515 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.034414
m1713 s72a net019535 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.077043
m1709 net015668 s71a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.025406
m1707 net019515 chal72 net015668 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.010213
m1705 vss! chal72 net019511 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.079686
m1704 net019515 net019511 net015683 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.022035
m1702 net015683 s71b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.021461
m1698 net019535 chal72 net015692 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.015506
m1697 net015692 s71b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.061221
m1695 net019535 net019531 net015699 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.034499
m1693 vss! chal72 net019531 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.033758
m1692 net015699 s71a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.018144
m1691 s71b net019563 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.014882
m1689 s71a net019583 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.142586
m1685 net015716 s70a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.061103
m1683 net019563 chal71 net015716 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.093795
m1681 vss! chal71 net019559 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.015080
m1680 net019563 net019559 net015731 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.062853
m1678 net015731 s70b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.004179
m1674 net019583 chal71 net015740 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.037395
m1673 net015740 s70b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.018144
m1671 net019583 net019579 net015747 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.067121
m1669 vss! chal71 net019579 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.088675
m1668 net015747 s70a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.067272
m1666 vss! chal70 net019599 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.039463
m1664 vss! chal70 net019603 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.090218
m1662 net015764 s69a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.028061
m1660 net019607 chal70 net015764 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.036959
m1658 s70b net019607 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.175879
m1657 net019607 net019599 net015779 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.001696
m1654 net015779 s69b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.146689
m1651 net019627 chal70 net015788 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.013191
m1650 net015788 s69b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.045093
m1648 net019627 net019603 net015795 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.070544
m1647 s70a net019627 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.126767
m1644 net015795 s69a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.034261
m1642 net015804 s68a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.021100
m1640 net019647 chal69 net015804 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.068874
m1638 net019647 net12759 net13288 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.017743
m1637 s69b net019647 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.055158
m1634 net13288 s68b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.041531
m1617 s68a net020396 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.034454
m1616 s68b net020408 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.039584
m1613 s67b net020444 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.002996
m1612 s67a net020456 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.136951
m1609 vss! chal68 net020380 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.089054
m1608 vss! chal68 net020384 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.019255
m1607 net017128 s67a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.064872
m1606 net020396 net020380 net017128 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.050523
m1605 net020396 chal68 net017133 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.030868
m1604 net017133 s67b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.076503
m1603 net017137 s67a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.011907
m1602 net020408 chal68 net017137 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.091339
m1601 net020408 net020384 net017148 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.065109
m1600 net017148 s67b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.023671
m1589 vss! chal67 net020420 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.037163
m1588 vss! chal67 net020424 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.053015
m1587 s66b net020484 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.184209
m1586 s66a net020496 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.053213
m1575 net017176 s66b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.131240
m1574 net020444 net020420 net017176 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.034975
m1573 net020444 chal67 net017181 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.096343
m1572 net017181 s66a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.004129
m1571 net017185 s66b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.086129
m1570 net020456 chal67 net017185 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.061073
m1569 net020456 net020424 net017196 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.056187
m1568 net017196 s66a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.077166
m1567 vss! chal66 net020468 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.033625
m1566 vss! chal66 net020472 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.006401
m1555 net017216 s65b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.093320
m1554 net020484 net020468 net017216 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.012815
m1553 net020484 chal66 net017221 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.113811
m1552 net017221 s65a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.049170
m1551 net017225 s65b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.053164
m1550 net020496 chal66 net017225 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.119676
m1549 net020496 net020472 net017236 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.033981
m1548 net017236 s65a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.006807
m1547 vss! chal65 net020508 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.075128
m1546 vss! chal65 net020512 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.050961
m1535 net017256 s64a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.171421
m1534 net020524 net020508 net017256 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.125410
m1533 net020524 chal65 net017261 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.058335
m1532 net017261 s64b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.061153
m1531 net017265 s64a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.112016
m1530 net020536 chal65 net017265 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.047478
m1529 net020536 net020512 net017276 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.065182
m1528 net017276 s64b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.077016
m1527 s65a net020524 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.042698
m1526 s65b net020536 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.089321
m1523 net017296 s63b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.029139
m1522 net020564 net020588 net017296 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.047948
m1521 net020564 chal64 net017301 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.018351
m1520 net017301 s63a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.016190
m1519 net017305 s63b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.103986
m1518 net020576 chal64 net017305 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.040623
m1517 net020576 net020592 net017316 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.025477
m1516 net017316 s63a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.042002
m1515 vss! chal64 net020588 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.059626
m1514 vss! chal64 net020592 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.055572
m1503 s64b net020564 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.007625
m1502 s64a net020576 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.108697
m1499 net017344 s62b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.151956
m1498 net020612 net020636 net017344 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.023919
m1497 net020612 chal63 net017349 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.018974
m1496 net017349 s62a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.024838
m1495 net017353 s62b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.091457
m1494 net020624 chal63 net017353 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.085480
m1493 net020624 net020640 net017364 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.017578
m1492 net017364 s62a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.010056
m1491 vss! chal63 net020636 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.094545
m1490 vss! chal63 net020640 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.011137
m1479 s63b net020612 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.120560
m1478 s63a net020624 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.001124
m1475 net017392 s61b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.081690
m1474 net020660 net020672 net017392 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.084884
m1473 net020660 chal62 net017397 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.018527
m1472 net017397 s61a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.118543
m1471 s62b net020660 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.076751
m1470 vss! chal62 net020672 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.004017
m1469 vss! chal62 net020676 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.013432
m1468 s62a net020688 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.089689
m1467 net017417 s61b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.028193
m1466 net020688 chal62 net017417 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.260555
m1465 net020688 net020676 net017428 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.116462
m1464 net017428 s61a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.057961
m1451 net017440 s60a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.090391
m1450 net16355 net020720 net017440 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.010742
m1449 net16355 chal61 net16352 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.010637
m1448 net16352 s60b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.048518
m1447 s61a net16355 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.081862
m1446 vss! chal61 net020720 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.055166
m1445 vss! chal61 net15733 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.024192
m1444 s61b net020736 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.046716
m1443 net017465 s60a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.062752
m1442 net020736 chal61 net017465 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.003823
m1441 net020736 net15733 net15780 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.097591
m1440 net15780 s60b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.021853
m1419 net017488 s59b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.058123
m1418 net020756 net020788 net017488 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.056965
m1417 net020756 chal60 net017493 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.136225
m1416 net017493 s59a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.028470
m1415 s60b net020756 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.032059
m1414 s60a net020768 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.031538
m1413 net017505 s59b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.012048
m1412 net020768 chal60 net017505 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.022126
m1411 net020768 net020792 net017516 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.000932
m1410 net017516 s59a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.042553
m1407 vss! chal60 net020788 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.050822
m1406 vss! chal60 net020792 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.052478
m1403 net017536 s58a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.092915
m1402 net020812 net020876 net017536 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.029334
m1401 net020812 chal59 net017541 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.071400
m1400 net017541 s58b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.023997
m1399 net017545 s58a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.027580
m1398 net020824 chal59 net017545 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.030977
m1397 net020824 net020880 net017556 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.053596
m1396 net017556 s58b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.145392
m1395 s59a net020812 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.007362
m1394 s59b net020824 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.002327
m1381 net017576 s57a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.019159
m1380 net020852 net020892 net017576 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.004880
m1379 net020852 chal58 net017581 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.022366
m1378 net017581 s57b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.073095
m1377 s58a net020852 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.034506
m1376 s58b net020864 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.100785
m1375 net017593 s57a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.012941
m1374 net020864 chal58 net017593 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.052090
m1373 net020864 net020896 net017604 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.003950
m1372 net017604 s57b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.071421
m1363 vss! chal59 net020876 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.124820
m1362 vss! chal59 net020880 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.098367
m1357 s57b net020916 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.007981
m1356 s57a net020928 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.030330
m1355 net017632 s56b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.038122
m1354 net020916 net020940 net017632 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.011824
m1353 net020916 chal57 net017637 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.041204
m1352 net017637 s56a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.126503
m1351 net017641 s56b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.084992
m1350 net020928 chal57 net017641 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.042448
m1349 net020928 net020944 net017652 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.019159
m1348 net017652 s56a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.082302
m1345 vss! chal58 net020892 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.041620
m1344 vss! chal58 net020896 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.026042
m1341 s56a net020972 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.063408
m1340 s56b net020984 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.016216
m1329 vss! chal57 net020940 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.005936
m1328 vss! chal57 net020944 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.042738
m1325 s55a net021012 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.058892
m1324 s55b net021024 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.114003
m1313 vss! chal56 net020956 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.033288
m1312 vss! chal56 net020960 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.021512
m1311 net017704 s55a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.016476
m1310 net020972 net020956 net017704 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.072383
m1309 net020972 chal56 net017709 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.023163
m1308 net017709 s55b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.035854
m1307 net017713 s55a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.037230
m1306 net020984 chal56 net017713 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.021454
m1305 net020984 net020960 net017724 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.062428
m1304 net017724 s55b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.102471
m1293 vss! chal55 net020996 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.092846
m1292 vss! chal55 net021000 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.051143
m1291 net017744 s54a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.016698
m1290 net021012 net020996 net017744 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.032752
m1289 net021012 chal55 net017749 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.049950
m1288 net017749 s54b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.099225
m1287 net017753 s54a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.074711
m1286 net021024 chal55 net017753 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.114267
m1285 net021024 net021000 net017764 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.068277
m1284 net017764 s54b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.048885
m1271 net017776 s53a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.004362
m1270 net021044 net021056 net017776 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.055909
m1269 net021044 chal54 net017781 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.010269
m1268 net017781 s53b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.082315
m1267 s54a net021044 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.004808
m1266 vss! chal54 net021056 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.120833
m1265 vss! chal54 net021060 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.101482
m1264 s54b net021072 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.019925
m1263 net017801 s53a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.061183
m1262 net021072 chal54 net017801 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.025795
m1261 net021072 net021060 net017812 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.088317
m1260 net017812 s53b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.123172
m1247 net14002 s52b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.027547
m1246 net021092 net13981 net14002 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.127053
m1245 net021092 chal53 net017829 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.062867
m1244 net017829 s52a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.038311
m1243 s53b net021092 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.116927
m1242 vss! chal53 net13981 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.039474
m1241 vss! chal53 net021108 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.021393
m1240 s53a net15177 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.043900
m1239 net15179 s52b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.097464
m1238 net15177 chal53 net15179 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.019271
m1237 net15177 net021108 net017860 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.011750
m1236 net017860 s52a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.152106
m1233 vss! chal52 net021132 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.091519
m1232 vss! chal52 net021136 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.030487
m1229 net017880 s51a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.122748
m1228 net021156 net021132 net017880 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.138466
m1227 net021156 chal52 net017885 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.010748
m1226 net017885 s51b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.103137
m1225 s52a net021156 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.064823
m1224 s52b net021168 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.018390
m1223 net017897 s51a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.100786
m1222 net021168 chal52 net017897 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.033148
m1221 net021168 net021136 net017908 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.007105
m1220 net017908 s51b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.029748
m1201 vss! chal51 net021212 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.014257
m1200 vss! chal51 net021216 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.049841
m1197 s51b net021188 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.017536
m1196 s51a net021200 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.013351
m1195 net017936 s50b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.155406
m1194 net021188 net021212 net017936 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.134274
m1193 net021188 chal51 net017941 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.074695
m1192 net017941 s50a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.005590
m1191 net017945 s50b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.014196
m1190 net021200 chal51 net017945 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.051179
m1189 net021200 net021216 net017956 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.091870
m1188 net017956 s50a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.079310
m1179 vss! chal50 net021260 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.012397
m1178 vss! chal50 net021264 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.232788
m1175 net017976 s49b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.025572
m1174 net021236 net021260 net017976 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.068837
m1173 net021236 chal50 net017981 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.004412
m1172 net017981 s49a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.120740
m1171 s50b net021236 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.131588
m1170 s50a net021248 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.074449
m1169 net017993 s49b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.005161
m1168 net021248 chal50 net017993 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.134457
m1167 net021248 net021264 net018004 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.044991
m1166 net018004 s49a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.025970
m1163 net018016 s48a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.010179
m1162 net021292 net021276 net018016 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.017164
m1161 net021292 chal49 net018021 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.132312
m1160 net018021 s48b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.032267
m1159 net018025 s48a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.015508
m1158 net021304 chal49 net018025 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.031890
m1157 net021304 net021280 net018036 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.028843
m1156 net018036 s48b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.012074
m1155 vss! chal49 net021276 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.043321
m1154 vss! chal49 net021280 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.006175
m1143 s49a net021292 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.053250
m1142 s49b net021304 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.115637
m1139 net018064 s47b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.060870
m1138 net021332 net021356 net018064 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.023131
m1137 net021332 chal48 net018069 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.005607
m1136 net018069 s47a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.117754
m1135 net018073 s47b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.070636
m1134 net021344 chal48 net018073 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.090556
m1133 net021344 net021360 net018084 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.186501
m1132 net018084 s47a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.149310
m1131 vss! chal48 net021356 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.051125
m1130 vss! chal48 net021360 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.058804
m1119 s48b net021332 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.001204
m1118 s48a net021344 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.069590
m1115 s47b net021388 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.002827
m1114 s47a net021400 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.028332
m1111 net018120 s46b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.079997
m1110 net021388 net021412 net018120 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.083867
m1109 net021388 chal47 net018125 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.083779
m1108 net018125 s46a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.006816
m1107 net018129 s46b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.043004
m1106 net021400 chal47 net018129 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.085302
m1105 net021400 net021416 net018140 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.040031
m1104 net018140 s46a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.008982
m1103 vss! chal47 net021412 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.112596
m1102 vss! chal47 net021416 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.066995
m1091 net018160 s45b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.140806
m1090 net021428 net021468 net018160 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.001406
m1089 net021428 chal46 net018165 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.031186
m1088 net018165 s45a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.101467
m1087 s46b net021428 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.077207
m1086 s46a net021448 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.061310
m1085 net018177 s45b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.064067
m1084 net021448 chal46 net018177 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.064038
m1083 net021448 net021472 net018188 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.075233
m1082 net018188 s45a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.009499
m1071 net018200 s44a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.031130
m1070 net14547 net021492 net018200 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.005776
m1069 net14547 chal45 net14549 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.072504
m1068 net14549 s44b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.011122
m1067 s45a net14547 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.021650
m1066 s45b net021504 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.162078
m1065 net018217 s44a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.046731
m1064 net021504 chal45 net018217 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.074661
m1063 net021504 net13381 net13404 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.044741
m1062 net13404 s44b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.053338
m1059 vss! chal46 net021468 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.029547
m1058 vss! chal46 net021472 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.034393
m1622 vss! chal69 net12759 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.046042
m1055 vss! chal45 net021492 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.100526
m1054 vss! chal45 net13381 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.107452
m1041 vss! chal44 net09677 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.122699
m1040 vss! chal44 net09681 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.089814
m1037 net07577 s43a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.006555
m1036 net09701 net09677 net07577 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.110607
m1035 net09701 chal44 net07582 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.017135
m1034 net07582 s43b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.071418
m1033 s44a net09701 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.078949
m1032 s44b net09713 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.156273
m1031 net07594 s43a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.054197
m1030 net09713 chal44 net07594 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.070102
m1029 net09713 net09681 net07605 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.079683
m1028 net07605 s43b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.001677
m1009 vss! chal43 net09757 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.095468
m1008 vss! chal43 net09761 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.086542
m1005 s43b net09733 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.010785
m1004 s43a net09745 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.055664
m1003 net07633 s42b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.040710
m1002 net09733 net09757 net07633 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.034836
m1001 net09733 chal43 net07638 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.065620
m1000 net07638 s42a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.080901
m999 net07642 s42b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.032846
m998 net09745 chal43 net07642 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.070309
m997 net09745 net09761 net07653 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.060189
m996 net07653 s42a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.023407
m987 vss! chal42 net09805 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.115743
m986 vss! chal42 net09809 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.048782
m983 net07673 s41b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.078555
m982 net09781 net09805 net07673 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.056445
m981 net09781 chal42 net07678 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.030350
m980 net07678 s41a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.028798
m979 s42b net09781 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.103591
m978 s42a net09793 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.093211
m977 net07690 s41b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.010689
m976 net09793 chal42 net07690 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.117411
m975 net09793 net09809 net07701 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.000600
m974 net07701 s41a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.124487
m971 net07713 s40a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.118305
m970 net09837 net09821 net07713 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.020397
m969 net09837 chal41 net07718 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.064708
m968 net07718 s40b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.050557
m967 net07722 s40a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.042828
m966 net09849 chal41 net07722 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.058449
m965 net09849 net09825 net07733 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.070916
m964 net07733 s40b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.034933
m963 vss! chal41 net09821 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.002857
m962 vss! chal41 net09825 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.010113
m951 s41a net09837 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.021164
m950 s41b net09849 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.051692
m947 net07761 s39b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.038530
m946 net09877 net09901 net07761 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.074513
m945 net09877 chal40 net07766 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.133376
m944 net07766 s39a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.011660
m943 net07770 s39b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.013841
m942 net09889 chal40 net07770 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.015452
m941 net09889 net09905 net07781 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.124099
m940 net07781 s39a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.086302
m939 vss! chal40 net09901 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.130466
m938 vss! chal40 net09905 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.015425
m927 s40b net09877 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.063604
m926 s40a net09889 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.041382
m923 s39b net09933 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.016169
m922 s39a net09945 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.122344
m919 net07817 s38b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.004888
m918 net09933 net09957 net07817 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.064889
m917 net09933 chal39 net07822 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.074072
m916 net07822 s38a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.015574
m915 net07826 s38b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.050686
m914 net09945 chal39 net07826 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.056589
m913 net09945 net09961 net07837 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.063168
m912 net07837 s38a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.004709
m911 vss! chal39 net09957 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.051772
m910 vss! chal39 net09961 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.027774
m899 net07857 s37b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.065505
m898 net09973 net09985 net07857 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.158004
m897 net09973 chal38 net07862 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.071549
m896 net07862 s37a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.012032
m895 s38b net09973 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.024354
m894 vss! chal38 net09985 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.080390
m893 vss! chal38 net09989 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.044774
m892 s38a net010001 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.042346
m891 net07882 s37b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.019961
m890 net010001 chal38 net07882 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.048665
m889 net010001 net09989 net07893 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.007450
m888 net07893 s37a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.078799
m875 net07905 s36a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.054035
m874 net6876 net010033 net07905 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.028779
m873 net6876 chal37 net6877 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.027103
m872 net6877 s36b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.115081
m871 s37a net6876 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.020747
m870 vss! chal37 net010033 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.121779
m869 vss! chal37 net5733 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.083845
m868 s37b net010049 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.044596
m867 net07930 s36a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.071173
m866 net010049 chal37 net07930 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.079035
m865 net010049 net5733 net5723 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.038956
m864 net5723 s36b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.052595
m1624 net015839 s68a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.115133
m843 net07953 s35b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.127579
m842 net010069 net010101 net07953 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.069815
m841 net010069 chal36 net07958 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.041531
m840 net07958 s35a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.019605
m839 s36b net010069 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.067695
m838 s36a net010081 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.004731
m837 net07970 s35b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.009793
m836 net010081 chal36 net07970 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.061242
m835 net010081 net010105 net07981 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.000665
m834 net07981 s35a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.077022
m831 net07993 s34a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.062349
m830 net010141 net010125 net07993 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.033406
m829 net010141 chal35 net07998 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.009711
m828 net07998 s34b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.112198
m827 net08002 s34a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.026427
m826 net010153 chal35 net08002 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.028430
m825 net010153 net010129 net08013 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.038030
m824 net08013 s34b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.084257
m823 vss! chal36 net010101 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.040629
m822 vss! chal36 net010105 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.004457
m821 s35a net010141 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.030313
m820 s35b net010153 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.041805
m813 net08041 s33a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.117846
m812 net010189 net010173 net08041 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.002921
m811 net010189 chal34 net08046 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.066027
m810 net08046 s33b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.015957
m809 s34a net010189 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.040377
m808 s34b net010201 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.012070
m807 net08058 s33a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.040952
m806 net010201 chal34 net08058 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.034543
m805 net010201 net010177 net08069 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.116988
m804 net08069 s33b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.027763
m803 vss! chal35 net010125 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.009871
m802 vss! chal35 net010129 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.083342
m787 s33b net010229 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.013520
m786 s33a net010241 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.101192
m785 vss! chal34 net010173 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.020201
m784 vss! chal34 net010177 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.086040
m763 s32a net010277 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.004478
m762 s32b net010289 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.010654
m761 vss! chal33 net010253 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.033918
m760 vss! chal33 net010257 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.114303
m759 net08121 s32b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.095823
m758 net010229 net010253 net08121 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.098973
m757 net010229 chal33 net08126 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.041351
m756 net08126 s32a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.054600
m755 net08130 s32b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.046007
m754 net010241 chal33 net08130 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.009227
m753 net010241 net010257 net08141 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.078569
m752 net08141 s32a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.016789
m741 vss! chal32 net010261 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.079951
m740 vss! chal32 net010265 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.077061
m739 net08161 s31a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.014622
m738 net010277 net010261 net08161 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.102626
m737 net010277 chal32 net08166 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.042440
m736 net08166 s31b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.086158
m735 net08170 s31a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.080042
m734 net010289 chal32 net08170 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.071797
m733 net010289 net010265 net08181 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.049632
m732 net08181 s31b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.007151
m721 vss! chal31 net010301 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.027659
m720 vss! chal31 net010305 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.036929
m719 net08201 s30a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.176717
m718 net010317 net010301 net08201 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.044567
m717 net010317 chal31 net08206 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.016410
m716 net08206 s30b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.048535
m715 net08210 s30a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.018517
m714 net010329 chal31 net08210 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.208498
m713 net010329 net010305 net08221 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.021092
m712 net08221 s30b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.055026
m709 s31a net010317 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.073162
m708 s31b net010329 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.022205
m695 net08241 s29a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.036436
m694 net010357 net010369 net08241 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.016659
m693 net010357 chal30 net08246 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.064531
m692 net08246 s29b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.137452
m691 s30a net010357 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.063800
m690 vss! chal30 net010369 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.146996
m689 vss! chal30 net010373 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.015012
m688 s30b net010385 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.055932
m687 net08266 s29a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.056724
m686 net010385 chal30 net08266 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.008244
m685 net010385 net010373 net08277 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.009662
m684 net08277 s29b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.028764
m1627 net13861 net019691 net015839 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.057890
m1620 vss! chal69 net019691 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.025312
m671 net5145 s28b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.071716
m670 net010405 net5123 net5145 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.048311
m669 net010405 chal29 net08294 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.053122
m668 net08294 s28a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.041332
m667 s29b net010405 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.024861
m666 vss! chal29 net5123 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.023850
m665 vss! chal29 net010421 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.015928
m664 s29a net6317 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.069919
m663 net6319 s28b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.022809
m662 net6317 chal29 net6319 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.041793
m661 net6317 net010421 net08325 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.009072
m660 net08325 s28a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.100824
m651 net08337 s27b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.057288
m650 net010453 net010485 net08337 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.020593
m649 net010453 chal28 net08342 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.080596
m648 net08342 s27a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.060219
m647 s28b net010453 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.003927
m646 s28a net010465 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.085032
m645 net08354 s27b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.065177
m644 net010465 chal28 net08354 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.101310
m643 net010465 net010489 net08365 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.065432
m642 net08365 s27a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.025734
m639 net08377 s26a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.016811
m638 net010525 net010509 net08377 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.040813
m637 net010525 chal27 net08382 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.071942
m636 net08382 s26b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.025379
m635 net08386 s26a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.054284
m634 net010537 chal27 net08386 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.052849
m633 net010537 net010513 net08397 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.165012
m632 net08397 s26b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.053004
m631 vss! chal28 net010485 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.104440
m630 vss! chal28 net010489 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.020704
m629 s27a net010525 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.046719
m628 s27b net010537 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.065986
m621 net08425 s25a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.057200
m620 net010573 net010557 net08425 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.034433
m619 net010573 chal26 net08430 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.001938
m618 net08430 s25b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.024164
m617 s26a net010573 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.015102
m616 s26b net010585 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.142030
m615 net08442 s25a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.112316
m614 net010585 chal26 net08442 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.059898
m613 net010585 net010561 net08453 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.083050
m612 net08453 s25b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.041342
m611 vss! chal27 net010509 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.034696
m610 vss! chal27 net010513 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.006230
m595 s25b net010613 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.072340
m594 s25a net010625 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.007047
m593 vss! chal26 net010557 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.116769
m592 vss! chal26 net010561 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.027940
m571 s24a net010661 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.043926
m570 s24b net010673 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.078494
m569 vss! chal25 net010637 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.064516
m568 vss! chal25 net010641 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.086733
m567 net08505 s24b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.100428
m566 net010613 net010637 net08505 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.065977
m565 net010613 chal25 net08510 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.062975
m564 net08510 s24a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.030944
m563 net08514 s24b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.115048
m562 net010625 chal25 net08514 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.035480
m561 net010625 net010641 net08525 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.054244
m560 net08525 s24a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.055561
m549 vss! chal24 net013341 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.022179
m548 vss! chal24 net010649 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.082024
m547 net08545 s23a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.000336
m546 net010661 net013341 net08545 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.029472
m545 net010661 chal24 net08550 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.110985
m544 net08550 s23b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.047922
m543 net08554 s23a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.009057
m542 net010673 chal24 net08554 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.076021
m541 net010673 net010649 net08565 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.156091
m540 net08565 s23b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.036188
m529 vss! chal23 net010685 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.059386
m528 vss! chal23 net013346 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.056980
m527 net08585 s22a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.087393
m526 net010701 net010685 net08585 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.047419
m525 net010701 chal23 net08590 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.005161
m524 net08590 s22b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.137321
m523 net08594 s22a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.111902
m522 net010713 chal23 net08594 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.003995
m521 net010713 net013346 net08605 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.042039
m520 net08605 s22b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.054982
m517 s23a net010701 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.030614
m516 s23b net010713 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.012586
m503 net08625 s21a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.037101
m502 net010741 net010753 net08625 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.174500
m501 net010741 chal22 net08630 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.138377
m500 net08630 s21b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.004157
m499 s22a net010741 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.099010
m498 vss! chal22 net010753 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.043441
m497 vss! chal22 net010757 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.024556
m496 s22b net010769 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.010110
m495 net08650 s21a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.053431
m494 net010769 chal22 net08650 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.085046
m493 net010769 net010757 net08661 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.043698
m492 net08661 s21b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.011804
m1628 s69a net13861 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.023013
m479 net3803 s20b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.072003
m478 net010789 net3767 net3803 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.027550
m477 net010789 chal21 net08678 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.108090
m476 net08678 s20a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.051370
m475 s21b net010789 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.067893
m474 vss! chal21 net3767 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.024474
m473 vss! chal21 net010805 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.011847
m472 s21a net4501 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.059357
m471 net4492 s20b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.074834
m470 net4501 chal21 net4492 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.020554
m469 net4501 net010805 net08709 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.076054
m468 net08709 s20a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.067292
m465 net09645 s19a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.111611
m464 net010633 net010617 net09645 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.051241
m463 net010633 chal20 net09650 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.011814
m462 net09650 s19b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.096699
m461 s20a net010633 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.065051
m460 s20b net010645 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.024419
m459 net09662 s19a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.018860
m458 net010645 chal20 net09662 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.035760
m457 net010645 net010621 net09673 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.172282
m456 net09673 s19b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.042979
m451 s19b net010665 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.027681
m450 s19a net010677 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.080133
m449 vss! chal20 net010617 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.156266
m448 vss! chal20 net010621 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.058803
m429 vss! chal19 net010689 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.042965
m428 vss! chal19 net010693 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.082051
m427 net09709 s18b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.067077
m426 net010665 net010689 net09709 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.066719
m425 net010665 chal19 net09714 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.049241
m424 net09714 s18a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.039193
m423 net09718 s18b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.072660
m422 net010677 chal19 net09718 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.012482
m421 net010677 net010693 net09729 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.032896
m420 net09729 s18a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.067192
m419 net3223 s17b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.031152
m418 net4091 net4123 net3223 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.113482
m417 net4091 chal18 net3228 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.011018
m416 net3228 s17a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.013822
m415 s18b net4091 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.058196
m414 s18a net4111 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.044613
m413 net3240 s17b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.073402
m412 net4111 chal18 net3240 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.017373
m411 net4111 net4127 net3251 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.036744
m410 net3251 s17a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.014926
m1630 net13861 chal69 net13857 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.167816
m399 vss! chal18 net4123 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.054069
m398 vss! chal18 net4127 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.028427
m397 net3271 s16a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.038732
m396 net4155 net4139 net3271 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.094708
m395 net4155 chal17 net3276 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.003018
m394 net3276 s16b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.011734
m393 s17a net4155 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.089572
m392 s17b net4167 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.007855
m391 net3288 s16a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.049384
m390 net4167 chal17 net3288 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.009128
m389 net4167 net4143 net3299 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.127783
m388 net3299 s16b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.103130
m383 vss! chal17 net4139 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.052598
m382 vss! chal17 net4143 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.030361
m381 s16b net4195 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.040345
m380 s16a net4207 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.058412
m367 net3327 s15b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.044016
m366 net4195 net4219 net3327 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.017910
m365 net4195 chal16 net3332 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.039343
m364 net3332 s15a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.085989
m363 net3336 s15b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.038783
m362 net4207 chal16 net3336 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.047619
m361 net4207 net4223 net3347 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.048382
m360 net3347 s15a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.015536
m359 vss! chal16 net4219 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.038215
m358 vss! chal16 net4223 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.032182
m357 s15b net4243 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.148170
m356 s15a net4255 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.007637
m343 net3375 s14b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.064388
m342 net4243 net4267 net3375 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.092652
m341 net4243 chal15 net3380 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.006906
m340 net3380 s14a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.028465
m339 net3384 s14b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.094632
m338 net4255 chal15 net3384 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.032887
m337 net4255 net4271 net3395 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.113961
m336 net3395 s14a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.047769
m335 vss! chal15 net4267 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.136060
m334 vss! chal15 net4271 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.051817
m323 net3415 s13b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.022622
m322 net4283 net4295 net3415 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.095175
m321 net4283 chal14 net3420 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.020372
m320 net3420 s13a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.155330
m319 s14b net4283 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.010124
m318 vss! chal14 net4295 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.005509
m317 vss! chal14 net4299 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.039355
m316 s14a net4311 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.011499
m315 net3440 s13b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.082159
m314 net4311 chal14 net3440 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.092988
m313 net4311 net4299 net3451 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.172145
m312 net3451 s13a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.094654
m299 net3463 s12a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.017274
m298 net4331 net4343 net3463 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.020161
m273 net4331 chal13 net3468 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.061087
m272 net3468 s12b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.065153
m271 s13a net4331 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.005331
m270 vss! chal13 net4343 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.068997
m269 vss! chal13 net4347 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.064809
m268 s13b net4359 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.149205
m267 net3488 s12a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.022808
m266 net4359 chal13 net3488 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.015611
m265 net4359 net4347 net3499 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.191401
m264 net3499 s12b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.021598
m1631 net13857 s68b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.010228
m11 net3511 start2 vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.002641
m10 net4379 net4391 net3511 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.045335
m9 net4379 chal1 net3516 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.090118
m8 net3516 start1 vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.028771
m7 s1b net4379 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.154038
m6 vss! chal1 net4391 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.065033
m_i_10 vss! chal1 net4395 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.000187
m_i_0 s1a net4407 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.081034
m_i_3 net3536 start2 vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.081517
m_i_2 net4407 chal1 net3536 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.055051
m_i_5 net4407 net4395 net3547 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.011224
m_i_4 net3547 start1 vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.003328
m12 net3559 s1a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.103521
m13 net4427 net4439 net3559 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.040444
m14 net4427 chal2 net3564 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.000247
m15 net3564 s1b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.009567
m16 s2a net4427 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.107729
m17 vss! chal2 net4439 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.034639
m18 vss! chal2 net4443 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.018820
m19 s2b net4455 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.039800
m20 net3584 s1a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.006901
m21 net4455 chal2 net3584 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.069106
m22 net4455 net4443 net3595 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.025733
m23 net3595 s1b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.113561
m36 vss! chal3 net4467 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.048590
m37 vss! chal3 net4471 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.074056
m40 net3615 s2a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.048620
m41 net4483 net4467 net3615 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.018908
m42 net4483 chal3 net3620 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.015069
m43 net3620 s2b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.019422
m44 s3a net4483 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.029652
m45 s3b net4503 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.035065
m46 net3632 s2a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.148720
m47 net4503 chal3 net3632 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.071481
m48 net4503 net4471 net3643 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.039054
m49 net3643 s2b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.019936
m60 vss! chal4 net4515 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.067870
m61 vss! chal4 net4519 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.075768
m64 net3663 s3a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.087932
m65 net4531 net4515 net3663 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.051882
m66 net4531 chal4 net3668 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.008567
m67 net3668 s3b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.025115
m68 s4a net4531 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.084364
m69 s4b net4551 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.031205
m70 net3680 s3a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.037263
m71 net4551 chal4 net3680 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.188502
m72 net4551 net4519 net3691 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.038825
m73 net3691 s3b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.082356
m94 net3703 s4b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.003548
m95 net4571 net4603 net3703 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.126159
m96 net4571 chal5 net3708 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.006657
m97 net3708 s4a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.069650
m98 s5b net4571 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.001165
m99 s5a net4591 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.120123
m100 net3720 s4b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.088032
m101 net4591 chal5 net3720 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.082891
m102 net4591 net4607 net3731 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.019715
m103 net3731 s4a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.064004
m106 vss! chal5 net4603 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.033792
m107 vss! chal5 net4607 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.026149
m108 vss! chal6 net4611 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.060513
m109 vss! chal6 net4615 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.003854
m112 net3759 s5a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.065128
m113 net4627 net4611 net3759 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.053451
m114 net4627 chal6 net3764 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.086499
m115 net3764 s5b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.048907
m116 s6a net4627 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.059811
m117 s6b net4647 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.019220
m118 net3776 s5a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.015601
m119 net4647 chal6 net3776 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.122138
m120 net4647 net4615 net3787 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.054084
m121 net3787 s5b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.048964
m142 net3799 s6b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.088615
m143 net4667 net4699 net3799 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.082178
m144 net4667 chal7 net3804 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.072793
m145 net3804 s6a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.109705
m146 s7b net4667 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.017491
m147 s7a net4687 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.067589
m148 net3816 s6b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.011602
m149 net4687 chal7 net3816 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.003198
m150 net4687 net4703 net3827 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.119669
m151 net3827 s6a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.025931
m154 vss! chal7 net4699 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.045952
m155 vss! chal7 net4703 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.058197
m166 net3847 s7b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.061320
m167 net4715 net4747 net3847 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.009682
m168 net4715 chal8 net3852 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.156956
m169 net3852 s7a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.011674
m170 s8b net4715 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.032133
m171 s8a net4735 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.038234
m172 net3864 s7b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.091161
m173 net4735 chal8 net3864 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.028807
m174 net4735 net4751 net3875 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.037805
m175 net3875 s7a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.095653
m178 vss! chal8 net4747 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.049479
m179 vss! chal8 net4751 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.042530
m180 vss! chal9 net4755 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.064387
m181 vss! chal9 net4759 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.062958
m184 net3903 s8a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.002290
m185 net4771 net4755 net3903 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.099110
m186 net4771 chal9 net3908 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.117660
m187 net3908 s8b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.002645
m188 net3912 s8a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.116442
m189 net4783 chal9 net3912 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.058170
m190 net4783 net4759 net3923 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.073336
m191 net3923 s8b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.125567
m200 s9a net4771 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.033959
m201 s9b net4783 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.044354
m204 vss! chal10 net4803 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.077133
m205 vss! chal10 net4807 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.050191
m216 net3951 s9a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.154002
m217 net4819 net4803 net3951 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.062343
m218 net4819 chal10 net3956 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.044480
m219 net3956 s9b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.026145
m220 s10a net4819 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.036531
m221 s10b net4831 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.049903
m222 net3968 s9a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.081788
m223 net4831 chal10 net3968 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.023798
m224 net4831 net4807 net3979 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.071031
m225 net3979 s9b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.006520
m228 vss! chal11 net4851 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.107534
m229 vss! chal11 net4855 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.040335
m232 net3999 s10a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.040044
m233 net4867 net4851 net3999 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.010268
m234 net4867 chal11 net4004 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.064801
m235 net4004 s10b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.089120
m236 s11a net4867 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.069154
m237 s11b net4887 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.049830
m238 net4016 s10a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.093401
m239 net4887 chal11 net4016 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.070297
m240 net4887 net4855 net4027 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.042596
m241 net4027 s10b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.002515
m286 net4032 s11b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.017875
m297 s12a net4915 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =0.048801
m296 s12b net4935 vss! vss! NMOS_VTL L=50e-9 W=415e-9 DELVTO =-0.030183
m285 net4044 s11a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.108774
m284 net4935 chal12 net4044 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.024266
m283 net4935 net4927 net4055 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.053654
m282 net4055 s11b vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.034542
m293 vss! chal12 net4923 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.105318
m292 vss! chal12 net4927 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.045490
m289 net4075 s11a vss! vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =-0.074234
m288 net4915 net4923 net4075 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.080831
m287 net4915 chal12 net4032 vss! NMOS_VTL L=50e-9 W=210e-9 DELVTO =0.022348
m3153 s128a net028885 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.154247
m3150 vdd! s127a net028294 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.018753
m3149 net028294 chal128 net028885 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.044664
m3146 s127a net028921 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.001356
m3142 vdd! s126a net028306 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.030258
m3141 net028306 chal127 net028921 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.111282
m3139 s126a net028965 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.017476
m3136 vdd! s125a net028318 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.053418
m3135 net028318 chal126 net028965 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.000401
m3130 s125a net21589 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.025178
m3128 net21858 chal125 net21589 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.001813
m3127 vdd! s124a net21858 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.146248
m3126 s124a net029037 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.086931
m3121 net028338 chal124 net029037 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.023950
m3120 vdd! s123a net028338 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.038541
m3119 s123a net029065 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.045829
m3117 vdd! s122a net028354 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.020077
m3116 net028354 chal123 net029065 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.099285
m3112 vdd! s121a net028362 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.078325
m3111 net028362 chal122 net029101 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.005228
m3107 s122a net029101 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.075888
m3102 s121a net029145 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.001018
m3100 net028374 chal121 net029145 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.045005
m3099 vdd! s120a net028374 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.113391
m3097 s120a net029173 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.024412
m3094 vdd! s119a net028390 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.075839
m3093 net028390 chal120 net029173 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.156808
m3090 s119a net029209 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.016495
m3086 vdd! s118a net028402 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.087722
m3085 net028402 chal119 net029209 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.072114
m3083 s118a net029245 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.041498
m3081 net028410 chal118 net029245 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.076318
m3079 vdd! s117a net028410 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.014662
m3075 s117a net20711 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.036345
m3072 net21789 chal117 net20711 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.126157
m3071 vdd! s116a net21789 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.006029
m3070 vdd! s115a net028434 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.026643
m3069 net028434 chal116 net029317 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.024355
m3065 s116a net029317 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.035513
m3060 s115a net029361 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.085552
m3058 net028446 chal115 net029361 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.001510
m3057 vdd! s114a net028446 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.062000
m3056 s114a net029389 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.013414
m3051 net028458 chal114 net029389 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.048266
m3050 vdd! s113a net028458 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.137153
m3049 s113a net029425 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.031643
m3047 vdd! s112a net028474 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.037328
m3046 net028474 chal113 net029425 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.031994
m3042 s112a net029469 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.006261
m3040 net028482 chal112 net029469 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.194781
m3039 vdd! s111a net028482 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.012693
m3035 net028490 chal111 net029497 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.041786
m3034 vdd! s110a net028490 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.070156
m3031 s111a net029497 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.064737
m3028 s110a net029533 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.106518
m3026 net028506 chal110 net029533 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.044806
m3025 vdd! s109a net028506 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.031361
m3021 s109a net19022 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.017757
m3020 vdd! s108a net21766 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.007344
m3019 net21766 chal109 net19022 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.039225
m3014 vdd! s107a net028530 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.030341
m3013 net028530 chal108 net029609 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.032953
m3009 s108a net029609 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.058980
m3006 s107a net029641 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.026314
m3004 net028542 chal107 net029641 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.078530
m3003 vdd! s106a net028542 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.057742
m3000 s106a net029677 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.014969
m2995 net028554 chal106 net029677 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.050402
m2994 vdd! s105a net028554 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.069543
m2993 s105a net029717 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.054731
m2989 vdd! s104a net028570 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.019339
m2988 net028570 chal105 net029717 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.005085
m2986 s104a net029749 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.019021
m2984 net028578 chal104 net029749 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.046987
m2983 vdd! s103a net028578 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.126190
m2979 net028586 chal103 net029785 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.062727
m2978 vdd! s102a net028586 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.002061
m2975 s103a net029785 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.052330
m2972 s102a net029821 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.005883
m2970 net028602 chal102 net029821 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.069833
m2969 vdd! s101a net028602 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.006115
m2965 s101a net19841 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.065945
m2964 vdd! s100a net20458 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.006125
m2963 net20458 chal101 net19841 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.083494
m2958 s100a net029893 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.034872
m2954 net028626 chal100 net029893 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.030628
m2953 vdd! s99a net028626 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.023103
m2951 s99a net029933 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.098010
m2947 vdd! s98a net028642 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.036532
m2946 net028642 chal99 net029933 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.070344
m2941 s98a net029965 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.079645
m2940 vdd! s97a net028654 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.010727
m2939 net028654 chal98 net029965 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.068197
m2936 s97a net030009 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.068565
m2933 net028662 chal97 net030009 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.064502
m2932 vdd! s96a net028662 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.057620
m2929 s96a net030045 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.000460
m2925 vdd! s95a net028678 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.026189
m2924 net028678 chal96 net030045 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.038864
m2922 s95a net030073 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.008725
m2919 vdd! s94a net028690 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.058588
m2918 net028690 chal95 net030073 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.090123
m2913 s94a net030109 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.053096
m2911 vdd! s93a net028702 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.071440
m2910 net028702 chal94 net030109 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.118610
m2908 s93a net20343 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.060423
m2905 net20337 chal93 net20343 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.030750
m2904 vdd! s92a net20337 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.087281
m2902 s92a net030181 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.046039
m2901 net028722 chal92 net030181 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.009319
m2900 vdd! s91a net028722 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.070965
m2895 s91a net030217 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.035628
m2891 net028734 chal91 net030217 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.088515
m2890 vdd! s90a net028734 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.011032
m2888 s90a net030261 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.062904
m2886 net028746 chal90 net030261 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.078258
m2885 vdd! s89a net028746 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.086932
m2881 s89a net030297 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.027892
m2876 net028758 chal89 net030297 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.023758
m2875 vdd! s88a net028758 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.054850
m2874 s88a net030325 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.052782
m2872 vdd! s87a net028774 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.074591
m2871 net028774 chal88 net030325 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.104115
m2867 s87a net030361 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.148941
m2863 vdd! s86a net028786 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.019164
m2862 net028786 chal87 net030361 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.052732
m2860 s86a net030397 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.000859
m2858 net028794 chal86 net030397 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.003435
m2857 vdd! s85a net028794 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.035596
m2853 s85a net030437 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.137568
m2849 vdd! s84a net028810 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.032223
m2848 net028810 chal85 net030437 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.048860
m2846 s84a net030469 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.084788
m2844 net028818 chal84 net030469 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.023783
m2843 vdd! s83a net028818 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.101405
m2839 s83a net030505 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.031074
m2835 net028830 chal83 net030505 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.104146
m2834 vdd! s82a net028830 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.032989
m2832 s82a net030541 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.010165
m2829 net028842 chal82 net030541 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.044655
m2828 vdd! s81a net028842 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.049890
m2825 s81a net19306 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.048794
m2821 net20133 chal81 net19306 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.101290
m2819 vdd! s80a net20133 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.106803
m2817 s128b net028869 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.094186
m2815 net028866 net028893 net028869 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.057641
m2812 net028870 chal128 net028869 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.028853
m2811 vdd! s127a net028866 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.108233
m2809 vdd! s127b net028870 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.129286
m2807 net028882 net028897 net028885 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.054061
m2805 vdd! s127b net028882 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.002933
m2804 vdd! chal128 net028893 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.030175
m2802 vdd! chal128 net028897 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.008426
m2797 s127b net028905 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.014196
m2793 net028902 net028929 net028905 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.013591
m2792 net028906 chal127 net028905 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.076060
m2791 vdd! s126a net028902 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.192411
m2790 vdd! s126b net028906 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.000412
m2789 net028918 net028933 net028921 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.017530
m2788 vdd! s126b net028918 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.032809
m2787 vdd! chal127 net028929 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.010081
m2785 vdd! chal127 net028933 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.037395
m2783 s126b net028949 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.019946
m2776 vdd! chal126 net028941 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.001269
m2774 vdd! chal126 net028945 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.115494
m2773 net028946 net028941 net028949 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.078000
m2772 vdd! s125a net028946 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.026132
m2771 net028954 chal126 net028949 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.011927
m2770 vdd! s125b net028954 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.074688
m2769 net028962 net028945 net028965 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.082645
m2768 vdd! s125b net028962 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.042904
m2766 s125b net028977 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.009438
m2764 net028974 net15878 net028977 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.096383
m2762 vdd! s124a net028974 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.038202
m2759 vdd! s124b net028986 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.081595
m2758 net028986 chal125 net028977 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.155300
m2756 net028990 net029005 net21589 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.009747
m2754 vdd! s124b net028990 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.015900
m2753 vdd! chal125 net15878 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.038819
m2751 vdd! chal125 net029005 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.063978
m2749 s124b net029021 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.014013
m2742 vdd! chal124 net029013 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.010415
m2741 vdd! s123a net029018 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.050495
m2740 net029018 net029013 net029021 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.084091
m2739 net029022 chal124 net029021 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.003632
m2737 vdd! s123b net029022 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.037281
m2736 vdd! chal124 net029033 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.032022
m2735 net029034 net029033 net029037 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.127279
m2734 vdd! s123b net029034 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.035557
m2732 s123b net029049 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.029431
m2731 net029046 net029073 net029049 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.023585
m2730 vdd! s122a net029046 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.031803
m2727 net029054 chal123 net029049 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.033058
m2725 vdd! s122b net029054 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.000446
m2723 net029062 net029077 net029065 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.119811
m2721 vdd! s122b net029062 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.016760
m2719 vdd! chal123 net029073 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.059041
m2717 vdd! chal123 net029077 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.028893
m2709 s122b net029085 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.082808
m2708 net029082 net029109 net029085 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.054706
m2707 net029086 chal122 net029085 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.082037
m2706 vdd! s121a net029082 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.014991
m2705 vdd! s121b net029086 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.010566
m2704 net029098 net029113 net029101 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.127002
m2703 vdd! s121b net029098 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.066192
m2702 vdd! chal122 net029109 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.007524
m2700 vdd! chal122 net029113 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.003923
m2698 s121b net029125 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.070945
m2691 vdd! chal121 net029121 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.019136
m2690 net029122 net029121 net029125 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.030159
m2689 vdd! s120a net029122 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.050249
m2687 vdd! s120b net029134 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.037229
m2686 net029134 chal121 net029125 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.037916
m2685 vdd! chal121 net029141 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.014824
m2684 net029142 net029141 net029145 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.109596
m2683 vdd! s120b net029142 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.037651
m2681 s120b net029157 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.203666
m2679 net029154 net029181 net029157 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.034498
m2677 vdd! s119a net029154 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.015057
m2674 net029162 chal120 net029157 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.028631
m2673 vdd! s119b net029162 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.127362
m2671 net029170 net029185 net029173 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.009492
m2669 vdd! s119b net029170 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.215527
m2668 vdd! chal120 net029181 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.064637
m2666 vdd! chal120 net029185 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.101859
m2664 s119b net029193 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.014931
m2662 net029190 net029217 net029193 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.075153
m2660 vdd! s118a net029190 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.036116
m2657 net029198 chal119 net029193 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.031057
m2656 vdd! s118b net029198 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.113858
m2654 net029206 net029221 net029209 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.037322
m2652 vdd! s118b net029206 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.082990
m2651 vdd! chal119 net029217 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.030064
m2649 vdd! chal119 net029221 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.040993
m2647 s118b net029229 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.099172
m2645 net029226 net029253 net029229 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.008216
m2643 vdd! s117a net029226 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.106320
m2640 net029234 chal118 net029229 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.005547
m2639 vdd! s117b net029234 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.050216
m2637 net029242 net029257 net029245 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.034716
m2635 vdd! s117b net029242 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.043242
m2634 vdd! chal118 net029253 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.023751
m2632 vdd! chal118 net029257 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.026911
m2626 s117b net029265 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.022858
m2623 net029262 net16859 net029265 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.008935
m2622 vdd! s116a net029262 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.009399
m2621 vdd! s116b net029274 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.008994
m2620 net029274 chal117 net029265 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.101901
m2619 net029278 net029293 net20711 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.001279
m2618 vdd! s116b net029278 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.083331
m2617 vdd! chal117 net16859 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.008956
m2615 vdd! chal117 net029293 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.081651
m2609 s116b net029301 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.095394
m2606 net029298 net029325 net029301 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.057468
m2605 vdd! s115a net029298 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.037744
m2604 net029306 chal116 net029301 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.144523
m2603 vdd! s115b net029306 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.079755
m2602 net029314 net029329 net029317 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.059738
m2601 vdd! s115b net029314 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.145093
m2600 vdd! chal116 net029325 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.088603
m2598 vdd! chal116 net029329 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.049160
m2596 s115b net029345 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.022939
m2589 vdd! chal115 net029337 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.091809
m2588 vdd! s114a net029342 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.045856
m2587 net029342 net029337 net029345 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.036590
m2586 net029346 chal115 net029345 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.011576
m2584 vdd! s114b net029346 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.038398
m2583 vdd! chal115 net029357 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.006178
m2582 net029358 net029357 net029361 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.096053
m2581 vdd! s114b net029358 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.128133
m2579 s114b net029377 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.067303
m2576 vdd! s113a net029374 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.032964
m2575 net029374 net029397 net029377 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.038832
m2573 net029378 chal114 net029377 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.071616
m2571 vdd! s113b net029378 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.036735
m2569 net029386 net029401 net029389 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.049244
m2567 vdd! s113b net029386 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.085955
m2566 vdd! chal114 net029397 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.073333
m2564 vdd! chal114 net029401 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.023953
m2559 s113b net029409 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.039894
m2555 net029406 net029433 net029409 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.001042
m2554 vdd! s112a net029406 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.069822
m2553 net029414 chal113 net029409 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.111967
m2552 vdd! s112b net029414 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.010737
m2551 net029422 net029437 net029425 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.050089
m2550 vdd! s112b net029422 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.050694
m2549 vdd! chal113 net029433 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.006023
m2547 vdd! chal113 net029437 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.115370
m2545 s112b net029453 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.012952
m2538 vdd! chal112 net029445 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.028209
m2537 vdd! s111a net029450 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.007366
m2536 net029450 net029445 net029453 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.043118
m2535 net029454 chal112 net029453 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.048127
m2534 vdd! s111b net029454 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.108973
m2532 vdd! chal112 net029465 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.072806
m2531 net029466 net029465 net029469 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.017378
m2530 vdd! s111b net029466 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.095256
m2528 s111b net029485 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.044567
m2527 vdd! s110a net029482 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.028213
m2526 net029482 net029505 net029485 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.005362
m2525 net029486 chal111 net029485 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.096771
m2524 vdd! s110b net029486 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.046260
m2523 net029494 net029509 net029497 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.100359
m2522 vdd! s110b net029494 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.044308
m2515 vdd! chal111 net029505 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.046803
m2513 vdd! chal111 net029509 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.122549
m2511 s110b net029517 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.005973
m2510 net029514 net029541 net029517 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.018411
m2508 vdd! s109a net029514 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.110279
m2507 net029522 chal110 net029517 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.032224
m2504 vdd! s109b net029522 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.104548
m2502 net029530 net029545 net029533 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.010358
m2500 vdd! s109b net029530 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.054563
m2498 vdd! chal110 net029541 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.090165
m2496 vdd! chal110 net029545 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.000314
m2494 s109b net029553 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.058849
m2493 net029550 net16774 net029553 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.088745
m2491 net029554 chal109 net029553 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.155917
m2490 vdd! s108a net029550 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.010686
m2487 vdd! s108b net029554 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.019758
m2485 net029566 net029581 net19022 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.137084
m2483 vdd! s108b net029566 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.104818
m2481 vdd! chal109 net16774 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.043668
m2479 vdd! chal109 net029581 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.027363
m2477 s108b net029589 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.014091
m2470 net029586 net029597 net029589 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.024049
m2469 vdd! s107a net029586 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.006047
m2468 vdd! chal108 net029597 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.009148
m2467 net029598 chal108 net029589 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.074484
m2466 vdd! s107b net029598 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.009289
m2464 net029606 net029613 net029609 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.104186
m2463 vdd! chal108 net029613 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.007600
m2462 vdd! s107b net029606 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.012781
m2460 s107b net029629 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.019491
m2459 vdd! s106a net029626 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.022800
m2458 net029626 net029649 net029629 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.061950
m2457 net029630 chal107 net029629 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.111580
m2456 vdd! s106b net029630 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.101875
m2455 net029638 net029653 net029641 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.043384
m2454 vdd! s106b net029638 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.029975
m2447 vdd! chal107 net029649 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.024199
m2445 vdd! chal107 net029653 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.024874
m2440 s106b net029665 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.040607
m2436 vdd! s105a net029662 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.145514
m2435 net029662 net029685 net029665 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.075533
m2434 net029666 chal106 net029665 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.059226
m2433 vdd! s105b net029666 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.128100
m2432 net029674 net029689 net029677 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.009353
m2431 vdd! s105b net029674 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.055636
m2430 vdd! chal106 net029685 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.026005
m2428 vdd! chal106 net029689 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.076303
m2426 s105b net029697 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.016209
m2419 net029694 net029705 net029697 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.017059
m2418 vdd! s104a net029694 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.070972
m2417 vdd! chal105 net029705 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.041154
m2416 net029706 chal105 net029697 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.022098
m2415 vdd! s104b net029706 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.099853
m2413 net029714 net029721 net029717 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.063984
m2412 vdd! chal105 net029721 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.032532
m2411 vdd! s104b net029714 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.020734
m2409 s104b net029737 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.024993
m2408 vdd! s103a net029734 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.039470
m2407 net029734 net029757 net029737 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.050427
m2404 net029738 chal104 net029737 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.035534
m2402 vdd! s103b net029738 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.027654
m2400 net029746 net029761 net029749 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.012836
m2398 vdd! s103b net029746 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.030506
m2396 vdd! chal104 net029757 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.032008
m2394 vdd! chal104 net029761 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.020377
m2392 s103b net029769 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.138159
m2391 net029766 net029793 net029769 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.023734
m2389 vdd! s102a net029766 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.075503
m2388 net029774 chal103 net029769 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.007833
m2385 vdd! s102b net029774 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.050223
m2383 net029782 net029797 net029785 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.000991
m2381 vdd! s102b net029782 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.087750
m2379 vdd! chal103 net029793 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.119123
m2377 vdd! chal103 net029797 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.055898
m2372 s102b net029805 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.111868
m2368 net029802 net029829 net029805 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.102704
m2367 vdd! s101a net029802 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.075255
m2366 net029810 chal102 net029805 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.017741
m2365 vdd! s101b net029810 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.170133
m2364 net029818 net029833 net029821 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.032267
m2363 vdd! s101b net029818 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.125558
m2362 vdd! chal102 net029829 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.077455
m2360 vdd! chal102 net029833 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.027806
m2358 s101b net029841 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.082079
m2351 net029838 net16703 net029841 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.039383
m2350 vdd! chal101 net16703 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.025476
m2349 net029846 chal101 net029841 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.045585
m2348 vdd! s100a net029838 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.098488
m2347 vdd! s100b net029846 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.188833
m2345 vdd! chal101 net029861 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.066753
m2344 net029862 net029861 net19841 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.100417
m2343 vdd! s100b net029862 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.046276
m2335 s100b net029881 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.075420
m2334 vdd! s99a net029878 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.140151
m2333 net029878 net029901 net029881 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.122317
m2332 net029882 chal100 net029881 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.033526
m2331 vdd! s99b net029882 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.066314
m2330 net029890 net029905 net029893 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.087724
m2329 vdd! s99b net029890 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.102933
m2328 vdd! chal100 net029901 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.027747
m2326 vdd! chal100 net029905 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.046033
m2324 s99b net029913 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.072363
m2317 net029910 net029921 net029913 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.038565
m2316 vdd! s98a net029910 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.053536
m2315 vdd! chal99 net029921 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.107110
m2314 net029922 chal99 net029913 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.009788
m2312 vdd! s98b net029922 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.037192
m2311 net029930 net029937 net029933 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.042151
m2310 vdd! chal99 net029937 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.080072
m2309 vdd! s98b net029930 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.083966
m2303 s98b net029949 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.034124
m2300 net029946 net029973 net029949 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.029310
m2299 vdd! s97a net029946 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.033436
m2298 net029954 chal98 net029949 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.082203
m2297 vdd! s97b net029954 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.081504
m2296 net029962 net029977 net029965 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.062885
m2295 vdd! s97b net029962 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.136314
m2294 vdd! chal98 net029973 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.057891
m2292 vdd! chal98 net029977 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.101574
m2286 s97b net029993 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.017698
m2283 vdd! chal97 net029985 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.025673
m2282 vdd! s96a net029990 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.014301
m2281 net029990 net029985 net029993 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.027191
m2280 net029994 chal97 net029993 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.030656
m2278 vdd! s96b net029994 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.012620
m2277 vdd! chal97 net030005 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.159910
m2276 net030006 net030005 net030009 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.074076
m2275 vdd! s96b net030006 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.173386
m2273 s96b net030029 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.066599
m2266 vdd! chal96 net030021 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.002274
m2264 vdd! chal96 net030025 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.034802
m2263 net030026 net030021 net030029 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.019933
m2262 vdd! s95a net030026 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.003211
m2261 net030034 chal96 net030029 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.022744
m2260 vdd! s95b net030034 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.092146
m2259 net030042 net030025 net030045 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.149083
m2258 vdd! s95b net030042 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.013729
m2256 s95b net030057 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.162726
m2253 net030054 net030081 net030057 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.062315
m2252 vdd! s94a net030054 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.018003
m2250 net030062 chal95 net030057 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.091619
m2248 vdd! s94b net030062 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.059892
m2246 net030070 net030085 net030073 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.063143
m2244 vdd! s94b net030070 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.052904
m2243 vdd! chal95 net030081 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.061283
m2241 vdd! chal95 net030085 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.010567
m2239 s94b net030093 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.030828
m2236 net030090 net030117 net030093 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.057935
m2235 vdd! s93a net030090 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.053853
m2233 net030098 chal94 net030093 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.108904
m2231 vdd! s93b net030098 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.108525
m2229 net030106 net030121 net030109 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.020352
m2227 vdd! s93b net030106 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.105912
m2226 vdd! chal94 net030117 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.050796
m2224 vdd! chal94 net030121 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.075293
m2216 s93b net030133 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.108417
m2215 vdd! s92a net030130 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.011376
m2214 net030130 net16587 net030133 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.022807
m2213 net030134 chal93 net030133 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.100934
m2212 vdd! s92b net030134 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.067205
m2211 net030142 net030157 net20343 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.024330
m2210 vdd! s92b net030142 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.007218
m2209 vdd! chal93 net16587 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.046244
m2207 vdd! chal93 net030157 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.080998
m2205 s92b net030169 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.064357
m2204 vdd! s91a net030166 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.067937
m2203 net030166 net030189 net030169 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.031927
m2200 net030170 chal92 net030169 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.008457
m2198 vdd! s91b net030170 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.000903
m2196 net030178 net030193 net030181 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.061989
m2194 vdd! s91b net030178 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.066401
m2192 vdd! chal92 net030189 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.031276
m2190 vdd! chal92 net030193 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.109210
m2185 s91b net030205 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.024256
m2181 vdd! s90a net030202 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.077572
m2180 net030202 net030225 net030205 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.095880
m2179 net030206 chal91 net030205 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.075040
m2178 vdd! s90b net030206 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.106149
m2177 net030214 net030229 net030217 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.025115
m2176 vdd! s90b net030214 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.112997
m2175 vdd! chal91 net030225 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.057664
m2173 vdd! chal91 net030229 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.010819
m2171 s90b net030245 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.101636
m2164 vdd! chal90 net030237 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.036694
m2163 vdd! s89a net030242 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.089229
m2162 net030242 net030237 net030245 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.054633
m2161 net030246 chal90 net030245 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.014209
m2160 vdd! s89b net030246 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.019690
m2158 vdd! chal90 net030257 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.129167
m2157 net030258 net030257 net030261 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.017628
m2156 vdd! s89b net030258 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.045175
m2154 s89b net030285 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.086194
m2147 vdd! chal89 net030273 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.061400
m2145 vdd! chal89 net030277 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.022858
m2144 vdd! s88a net030282 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.036705
m2143 net030282 net030273 net030285 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.033052
m2142 net030286 chal89 net030285 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.019231
m2141 vdd! s88b net030286 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.047091
m2140 net030294 net030277 net030297 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.040197
m2139 vdd! s88b net030294 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.049164
m2137 s88b net030309 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.017591
m2136 net030306 net030333 net030309 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.024669
m2135 vdd! s87a net030306 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.100302
m2132 net030314 chal88 net030309 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.077662
m2130 vdd! s87b net030314 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.014963
m2128 net18777 net030337 net030325 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.120848
m2126 vdd! s87b net18777 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.008878
m2124 vdd! chal88 net030333 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.054902
m2122 vdd! chal88 net030337 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.074703
m2120 s87b net030345 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.014360
m2119 net030342 net030369 net030345 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.086003
m2117 net030346 chal87 net030345 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.115905
m2116 vdd! s86a net030342 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.000143
m2113 vdd! s86b net030346 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.104008
m2111 net030358 net030373 net030361 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.011099
m2109 vdd! s86b net030358 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.061175
m2107 vdd! chal87 net030369 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.007269
m2105 vdd! chal87 net030373 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.121982
m2097 s86b net030381 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.057838
m2096 net030378 net030405 net030381 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.043486
m2095 vdd! s85a net030378 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.096490
m2094 net030386 chal86 net030381 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.015579
m2093 vdd! s85b net030386 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.143090
m2092 net030394 net030409 net030397 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.031159
m2091 vdd! s85b net030394 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.024755
m2090 vdd! chal86 net030405 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.015661
m2088 vdd! chal86 net030409 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.062408
m2086 s85b net030417 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.011863
m2079 net030414 net030421 net030417 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.026330
m2078 vdd! chal85 net030421 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.109008
m2077 net030422 chal85 net030417 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.036046
m2076 vdd! s84a net030414 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.011549
m2075 vdd! s84b net030422 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.018340
m2073 net030434 net030441 net030437 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.036428
m2072 vdd! chal85 net030441 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.047978
m2071 vdd! s84b net030434 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.041898
m2070 s84b net030453 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.024905
m2068 net030450 net030477 net030453 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.046773
m2066 vdd! s83a net030450 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.008775
m2064 vdd! s83b net030462 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.064426
m2063 net030462 chal84 net030453 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.016705
m2060 net030466 net030481 net030469 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.075404
m2058 vdd! s83b net030466 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.152463
m2056 vdd! chal84 net030477 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.007980
m2054 vdd! chal84 net030481 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.009880
m2053 s83b net030489 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.024497
m2051 net030486 net030513 net030489 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.026507
m2049 vdd! s82a net030486 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.023673
m2047 vdd! s82b net030498 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.038786
m2046 net030498 chal83 net030489 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.017871
m2043 net030502 net030517 net030505 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.080370
m2041 vdd! s82b net030502 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.006354
m2039 vdd! chal83 net030513 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.075546
m2037 vdd! chal83 net030517 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.007236
m2036 s82b net030525 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.030387
m2034 net030522 net030549 net030525 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.018916
m2032 vdd! s81a net030522 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.116290
m2030 vdd! s81b net030534 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.030882
m2029 net030534 chal82 net030525 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.029755
m2026 net030538 net030553 net030541 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.114077
m2024 vdd! s81b net030538 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.020905
m2022 vdd! chal82 net030549 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.037472
m2020 vdd! chal82 net030553 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.093354
m2017 s81b net030561 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.045863
m2011 net030558 net15612 net030561 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.012999
m2010 vdd! s80a net030558 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.060864
m2009 net030566 chal81 net030561 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.055766
m2008 vdd! s80b net030566 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.016720
m2007 net030574 net030589 net19306 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.081439
m2006 vdd! s80b net030574 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.035652
m2005 vdd! chal81 net15612 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.156496
m2003 vdd! chal81 net030589 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.011378
m1907 net019116 net019159 net019119 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.028159
m1905 vdd! s79a net019116 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.116276
m1903 s80b net019119 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.065660
m1902 vdd! s79b net019132 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.026361
m1901 net019132 chal80 net019119 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.002295
m1897 net019136 net019163 net019139 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.042490
m1896 vdd! s79b net019136 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.076233
m1893 net019144 chal80 net019139 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.067744
m1890 s80a net019139 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.021311
m1889 vdd! s79a net019144 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.013240
m1887 vdd! chal80 net019159 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.117320
m1885 vdd! chal80 net019163 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.120652
m1881 s79b net019179 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.121249
m1873 s79a net019199 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.001387
m1871 vdd! chal79 net019175 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.031719
m1870 net019176 net019175 net019179 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.046695
m1869 vdd! s78a net019176 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.074339
m1868 vdd! s78b net019188 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.140759
m1867 net019188 chal79 net019179 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.041456
m1865 vdd! chal79 net019195 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.005894
m1864 net019196 net019195 net019199 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.001242
m1863 vdd! s78b net019196 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.028427
m1862 net019204 chal79 net019199 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.021809
m1860 vdd! s78a net019204 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.133123
m1859 s78b net019227 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.010769
m1856 s78a net019247 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.035755
m1855 vdd! chal78 net019223 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.151991
m1854 net019224 net019223 net019227 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.104114
m1852 vdd! s77a net019224 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.054719
m1850 vdd! s77b net019236 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.010275
m1849 net019236 chal78 net019227 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.025316
m1845 vdd! chal78 net019243 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.175685
m1844 net019244 net019243 net019247 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.123013
m1843 vdd! s77b net019244 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.120970
m1840 net019252 chal78 net019247 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.019683
m1837 vdd! s77a net019252 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.060860
m1835 s77b net019279 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.072701
m1832 s77a net019295 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.066703
m1831 vdd! chal77 net019271 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.029867
m1829 vdd! chal77 net019275 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.032797
m1827 net019276 net019271 net019279 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.014241
m1825 vdd! s76a net019276 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.112046
m1823 vdd! s76b net019288 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.053610
m1822 net019288 chal77 net019279 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.017941
m1819 net019292 net019275 net019295 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.046351
m1818 vdd! s76b net019292 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.010723
m1815 net019300 chal77 net019295 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.027534
m1813 vdd! s76a net019300 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.077347
m1811 net019308 net019315 net019311 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.007146
m1810 vdd! chal76 net019315 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.120728
m1808 vdd! s75a net019308 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.058403
m1806 net019320 chal76 net019311 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.038253
m1805 s76b net019311 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.129164
m1801 vdd! s75b net019320 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.042702
m1799 vdd! s75b net13983 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.045790
m1798 net13983 net019343 net019339 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.023872
m1797 vdd! chal76 net019343 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.059028
m1794 net019344 chal76 net019339 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.051093
m1790 s76a net019339 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.090763
m1789 vdd! s75a net019344 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.057657
m1787 net019356 net019399 net019359 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.082735
m1785 vdd! s74a net019356 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.041878
m1783 net019364 chal75 net019359 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.004170
m1782 s75b net019359 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.109017
m1779 vdd! s74b net019364 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.034910
m1777 vdd! s74b net019380 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.014101
m1776 net019380 net019403 net019383 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.048394
m1773 net019384 chal75 net019383 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.013959
m1770 s75a net019383 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.032382
m1769 vdd! s74a net019384 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.026485
m1767 vdd! chal75 net019399 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.012383
m1765 vdd! chal75 net019403 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.113393
m1763 net019404 net019447 net019407 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.141504
m1761 vdd! s73a net019404 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.002405
m1759 net019412 chal74 net019407 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.054184
m1757 vdd! s73b net019412 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.006358
m1755 net019420 net019451 net019423 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.040420
m1754 vdd! s73b net019420 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.050299
m1751 net019428 chal74 net019423 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.138207
m1749 vdd! s73a net019428 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.108506
m1746 s74b net019407 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.002056
m1744 s74a net019423 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.045296
m1743 vdd! chal74 net019447 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.092560
m1741 vdd! chal74 net019451 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.129584
m1735 s73b net019463 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.065008
m1729 s73a net019487 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.035193
m1727 net019460 net019467 net019463 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.032830
m1726 vdd! chal73 net019467 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.030815
m1725 vdd! s72a net019460 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.070240
m1724 net019472 chal73 net019463 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.165987
m1722 vdd! s72b net019472 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.033308
m1721 vdd! s72b net019484 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.032868
m1720 net019484 net019491 net019487 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.008468
m1719 vdd! chal73 net019491 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.095844
m1718 net019492 chal73 net019487 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.066903
m1717 vdd! s72a net019492 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.051588
m1714 s72b net019515 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.013326
m1712 s72a net019535 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.005754
m1711 vdd! chal72 net019511 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.005155
m1710 net019512 net019511 net019515 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.012487
m1708 vdd! s71a net019512 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.054029
m1706 net019520 chal72 net019515 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.025223
m1703 vdd! s71b net019520 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.111229
m1701 vdd! chal72 net019531 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.080132
m1700 net019532 net019531 net019535 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.022537
m1699 vdd! s71b net019532 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.056061
m1696 net019540 chal72 net019535 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.046602
m1694 vdd! s71a net019540 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.115636
m1690 s71b net019563 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.081602
m1688 s71a net019583 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.005340
m1687 vdd! chal71 net019559 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.008884
m1686 net019560 net019559 net019563 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.006735
m1684 vdd! s70a net019560 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.049753
m1682 net019568 chal71 net019563 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.025897
m1679 vdd! s70b net019568 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.062816
m1677 vdd! chal71 net019579 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.004660
m1676 net019580 net019579 net019583 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.035772
m1675 vdd! s70b net019580 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.045876
m1672 net019588 chal71 net019583 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.071971
m1670 vdd! s70a net019588 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.037448
m1667 vdd! chal70 net019599 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.052168
m1665 vdd! chal70 net019603 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.026561
m1663 net019604 net019599 net019607 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.065998
m1661 vdd! s69a net019604 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.082292
m1659 net019612 chal70 net019607 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.075134
m1656 s70b net019607 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.076413
m1655 vdd! s69b net019612 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.113851
m1653 net019624 net019603 net019627 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.090195
m1652 vdd! s69b net019624 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.082748
m1649 net019632 chal70 net019627 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.036329
m1646 vdd! s69a net019632 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.008096
m1645 s70a net019627 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.016658
m1643 net019644 net12759 net019647 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.012999
m1641 vdd! s68a net019644 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.061804
m1639 net019652 chal69 net019647 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.045269
m1636 vdd! s68b net019652 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.042686
m1635 s69b net019647 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.216322
m1619 s68a net020396 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.111405
m1618 s68b net020408 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.076108
m1615 s67b net020444 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.067061
m1614 s67a net020456 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.001776
m1611 vdd! chal68 net020380 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.121769
m1610 vdd! chal68 net020384 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.013372
m1599 net020385 chal68 net020396 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.053301
m1598 vdd! s67a net020385 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.047009
m1597 net020393 net020380 net020396 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.112310
m1596 vdd! s67b net020393 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.085551
m1595 vdd! s67a net020405 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.031768
m1594 net020405 net020384 net020408 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.038621
m1593 vdd! s67b net020413 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.019787
m1592 net020413 chal68 net020408 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.035743
m1591 vdd! chal67 net020420 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.032971
m1590 vdd! chal67 net020424 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.031133
m1585 s66b net020484 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.101806
m1584 s66a net020496 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.009365
m1583 net020433 chal67 net020444 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.110687
m1582 vdd! s66b net020433 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.153493
m1581 net020441 net020420 net020444 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.017164
m1580 vdd! s66a net020441 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.033534
m1579 vdd! s66b net020453 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.027819
m1578 net020453 net020424 net020456 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.009773
m1577 vdd! s66a net020461 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.002606
m1576 net020461 chal67 net020456 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.071337
m1565 vdd! chal66 net020468 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.001774
m1564 vdd! chal66 net020472 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.153696
m1563 net020473 chal66 net020484 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.065371
m1562 vdd! s65b net020473 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.027592
m1561 net020481 net020468 net020484 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.019417
m1560 vdd! s65a net020481 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.019447
m1559 vdd! s65b net020493 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.088673
m1558 net020493 net020472 net020496 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.117763
m1557 vdd! s65a net020501 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.031147
m1556 net020501 chal66 net020496 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.057860
m1545 vdd! chal65 net020508 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.037328
m1544 vdd! chal65 net020512 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.087688
m1543 net020513 chal65 net020524 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.078978
m1542 vdd! s64a net020513 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.007174
m1541 net020521 net020508 net020524 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.101892
m1540 vdd! s64b net020521 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.090210
m1539 vdd! s64a net020533 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.025627
m1538 net020533 net020512 net020536 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.036443
m1537 vdd! s64b net020541 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.041259
m1536 net020541 chal65 net020536 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.109818
m1525 s65a net020524 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.092469
m1524 s65b net020536 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.031679
m1513 net020553 chal64 net020564 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.070026
m1512 vdd! s63b net020553 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.030597
m1511 net020561 net020588 net020564 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.091368
m1510 vdd! s63a net020561 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.003860
m1509 vdd! s63b net020573 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.047171
m1508 net020573 net020592 net020576 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.048001
m1507 vdd! s63a net020581 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.048602
m1506 net020581 chal64 net020576 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.022423
m1505 vdd! chal64 net020588 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.072649
m1504 vdd! chal64 net020592 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.047718
m1501 s64b net020564 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.092807
m1500 s64a net020576 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.024068
m1489 net020601 chal63 net020612 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.031826
m1488 vdd! s62b net020601 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.034217
m1487 net020609 net020636 net020612 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.108056
m1486 vdd! s62a net020609 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.033491
m1485 vdd! s62b net020621 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.039307
m1484 net020621 net020640 net020624 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.014076
m1483 vdd! s62a net020629 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.035213
m1482 net020629 chal63 net020624 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.070727
m1481 vdd! chal63 net020636 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.143906
m1480 vdd! chal63 net020640 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.027229
m1477 s63b net020612 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.037256
m1476 s63a net020624 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.067522
m1463 net020649 chal62 net020660 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.004777
m1462 vdd! s61b net020649 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.114230
m1461 net020657 net020672 net020660 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.028596
m1460 vdd! s61a net020657 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.022226
m1459 s62b net020660 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.033268
m1458 vdd! chal62 net020672 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.073744
m1457 vdd! chal62 net020676 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.084555
m1456 s62a net020688 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.185503
m1455 vdd! s61b net020685 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.013329
m1454 net020685 net020676 net020688 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.017424
m1453 vdd! s61a net020693 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.106623
m1452 net020693 chal62 net020688 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.018249
m1439 net16326 chal61 net16355 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.006427
m1438 vdd! s60a net16326 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.046933
m1437 net020705 net020720 net16355 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.043293
m1436 vdd! s60b net020705 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.070980
m1435 s61a net16355 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.016094
m1434 vdd! chal61 net020720 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.124365
m1433 vdd! chal61 net15733 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.035388
m1432 s61b net020736 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.072545
m1431 vdd! s60a net020733 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.108893
m1430 net020733 net15733 net020736 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.004098
m1429 vdd! s60b net020741 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.033488
m1428 net020741 chal61 net020736 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.016417
m1427 net020745 chal60 net020756 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.037163
m1426 vdd! s59b net020745 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.052793
m1425 net020753 net020788 net020756 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.047731
m1424 vdd! s59a net020753 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.014554
m1423 vdd! s59b net020765 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.018574
m1422 net020765 net020792 net020768 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.038659
m1421 vdd! s59a net020773 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.105679
m1420 net020773 chal60 net020768 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.050398
m1409 s60b net020756 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.080679
m1408 s60a net020768 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.043832
m1405 vdd! chal60 net020788 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.048598
m1404 vdd! chal60 net020792 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.089498
m1393 s59a net020812 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.089386
m1392 s59b net020824 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.121054
m1391 net020801 chal59 net020812 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.004699
m1390 vdd! s58a net020801 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.064664
m1389 net020809 net020876 net020812 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.074698
m1388 vdd! s58b net020809 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.067091
m1387 vdd! s58a net020821 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.107397
m1386 net020821 net020880 net020824 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.020414
m1385 vdd! s58b net020829 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.053806
m1384 net020829 chal59 net020824 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.092421
m1383 s58a net020852 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.039039
m1382 s58b net020864 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.000626
m1371 net020841 chal58 net020852 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.050901
m1370 vdd! s57a net020841 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.020327
m1369 net020849 net020892 net020852 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.044733
m1368 vdd! s57b net020849 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.147440
m1367 vdd! s57a net020861 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.054747
m1366 net020861 net020896 net020864 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.047775
m1365 vdd! s57b net020869 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.075349
m1364 net020869 chal58 net020864 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.017194
m1361 vdd! chal59 net020876 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.064898
m1360 vdd! chal59 net020880 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.022597
m1359 s57b net020916 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.101658
m1358 s57a net020928 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.104939
m1347 vdd! chal58 net020892 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.040832
m1346 vdd! chal58 net020896 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.001411
m1343 s56a net020972 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.042089
m1342 s56b net020984 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.089833
m1339 net020905 chal57 net020916 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.010336
m1338 vdd! s56b net020905 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.036038
m1337 net020913 net020940 net020916 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.002093
m1336 vdd! s56a net020913 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.093308
m1335 vdd! s56b net020925 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.037254
m1334 net020925 net020944 net020928 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.060167
m1333 vdd! s56a net020933 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.012761
m1332 net020933 chal57 net020928 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.017089
m1331 vdd! chal57 net020940 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.080196
m1330 vdd! chal57 net020944 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.013750
m1327 s55a net021012 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.079347
m1326 s55b net021024 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.030748
m1323 vdd! chal56 net020956 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.069665
m1322 vdd! chal56 net020960 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.014512
m1321 net020961 chal56 net020972 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.171168
m1320 vdd! s55a net020961 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.030635
m1319 net020969 net020956 net020972 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.014117
m1318 vdd! s55b net020969 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.080207
m1317 vdd! s55a net020981 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.071056
m1316 net020981 net020960 net020984 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.087803
m1315 vdd! s55b net020989 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.028058
m1314 net020989 chal56 net020984 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.058289
m1303 vdd! chal55 net020996 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.037366
m1302 vdd! chal55 net021000 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.121150
m1301 net021001 chal55 net021012 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.083524
m1300 vdd! s54a net021001 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.048029
m1299 net021009 net020996 net021012 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.128045
m1298 vdd! s54b net021009 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.019561
m1297 vdd! s54a net021021 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.056463
m1296 net021021 net021000 net021024 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.012451
m1295 vdd! s54b net021029 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.000341
m1294 net021029 chal55 net021024 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.142170
m1283 net021033 chal54 net021044 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.107703
m1282 vdd! s53a net021033 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.106221
m1281 net021041 net021056 net021044 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.056832
m1280 vdd! s53b net021041 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.151449
m1279 s54a net021044 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.057516
m1278 vdd! chal54 net021056 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.091491
m1277 vdd! chal54 net021060 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.104048
m1276 s54b net021072 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.002277
m1275 vdd! s53a net021069 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.041913
m1274 net021069 net021060 net021072 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.065288
m1273 vdd! s53b net021077 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.044329
m1272 net021077 chal54 net021072 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.056265
m1259 net021081 chal53 net021092 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.053501
m1258 vdd! s52b net021081 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.075418
m1257 net021089 net13981 net021092 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.026097
m1256 vdd! s52a net021089 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.083012
m1255 s53b net021092 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.080577
m1254 vdd! chal53 net13981 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.003965
m1253 vdd! chal53 net021108 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.138463
m1252 s53a net15177 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.064102
m1251 vdd! s52b net021117 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.103352
m1250 net021117 net021108 net15177 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.046294
m1249 vdd! s52a net15147 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.080323
m1248 net15147 chal53 net15177 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.016834
m1235 vdd! chal52 net021132 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.156639
m1234 vdd! chal52 net021136 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.088038
m1231 s52a net021156 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.038206
m1230 s52b net021168 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.061188
m1219 net021145 chal52 net021156 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.094039
m1218 vdd! s51a net021145 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.013445
m1217 net021153 net021132 net021156 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.007456
m1216 vdd! s51b net021153 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.018884
m1215 vdd! s51a net021165 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.011307
m1214 net021165 net021136 net021168 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.016259
m1213 vdd! s51b net021173 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.053488
m1212 net021173 chal52 net021168 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.065076
m1211 net021177 chal51 net021188 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.042551
m1210 vdd! s50b net021177 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.039558
m1209 net021185 net021212 net021188 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.065883
m1208 vdd! s50a net021185 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.095994
m1207 vdd! s50b net021197 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.096150
m1206 net021197 net021216 net021200 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.048063
m1205 vdd! s50a net021205 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.025484
m1204 net021205 chal51 net021200 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.043334
m1203 vdd! chal51 net021212 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.085078
m1202 vdd! chal51 net021216 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.018678
m1199 s51b net021188 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.050782
m1198 s51a net021200 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.202717
m1187 net021225 chal50 net021236 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.023476
m1186 vdd! s49b net021225 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.031333
m1185 net021233 net021260 net021236 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.021383
m1184 vdd! s49a net021233 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.078186
m1183 vdd! s49b net021245 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.028016
m1182 net021245 net021264 net021248 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.029201
m1181 vdd! s49a net021253 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.046409
m1180 net021253 chal50 net021248 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.001523
m1177 vdd! chal50 net021260 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.047925
m1176 vdd! chal50 net021264 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.151677
m1165 s50b net021236 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.098551
m1164 s50a net021248 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.037846
m1153 vdd! chal49 net021276 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.055182
m1152 vdd! chal49 net021280 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.048925
m1151 net021281 chal49 net021292 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.038233
m1150 vdd! s48a net021281 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.071948
m1149 net021289 net021276 net021292 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.013956
m1148 vdd! s48b net021289 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.026710
m1147 vdd! s48a net021301 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.004330
m1146 net021301 net021280 net021304 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.031446
m1145 vdd! s48b net021309 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.012985
m1144 net021309 chal49 net021304 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.072294
m1141 s49a net021292 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.109318
m1140 s49b net021304 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.165335
m1129 net021321 chal48 net021332 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.018918
m1128 vdd! s47b net021321 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.086247
m1127 net021329 net021356 net021332 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.080152
m1126 vdd! s47a net021329 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.002889
m1125 vdd! s47b net021341 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.091126
m1124 net021341 net021360 net021344 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.066031
m1123 vdd! s47a net021349 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.029332
m1122 net021349 chal48 net021344 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.057804
m1121 vdd! chal48 net021356 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.066827
m1120 vdd! chal48 net021360 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.038617
m1117 s48b net021332 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.055826
m1116 s48a net021344 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.152348
m1113 s47b net021388 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.019563
m1112 s47a net021400 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.091574
m1101 net021377 chal47 net021388 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.067024
m1100 vdd! s46b net021377 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.014719
m1099 net021385 net021412 net021388 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.094738
m1098 vdd! s46a net021385 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.007986
m1097 vdd! s46b net021397 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.038224
m1096 net021397 net021416 net021400 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.108764
m1095 vdd! s46a net021405 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.085537
m1094 net021405 chal47 net021400 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.053566
m1093 vdd! chal47 net021412 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.024787
m1092 vdd! chal47 net021416 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.028712
m1081 net021417 chal46 net021428 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.026897
m1080 vdd! s45b net021417 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.184034
m1079 net021425 net021468 net021428 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.025221
m1078 vdd! s45a net021425 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.075591
m1077 s46b net021428 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.033063
m1076 s46a net021448 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.002138
m1075 vdd! s45b net021445 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.107240
m1074 net021445 net021472 net021448 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.006954
m1073 vdd! s45a net021453 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.015805
m1072 net021453 chal46 net021448 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.036704
m1061 s45a net14547 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.043799
m1060 s45b net021504 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.094464
m1057 vdd! chal46 net021468 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.005290
m1056 vdd! chal46 net021472 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.035091
m1621 vdd! chal69 net019691 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.025263
m1053 net14553 chal45 net14547 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.046242
m1052 vdd! s44a net14553 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.065572
m1051 net021481 net021492 net14547 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.059634
m1050 vdd! s44b net021481 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.046839
m1049 vdd! chal45 net021492 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.043208
m1048 vdd! chal45 net13381 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.019855
m1047 vdd! s44a net021501 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.024568
m1046 net021501 net13381 net021504 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.071225
m1045 vdd! s44b net021509 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.047436
m1044 net021509 chal45 net021504 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.012191
m1043 vdd! chal44 net09677 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.011312
m1042 vdd! chal44 net09681 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.155966
m1039 s44a net09701 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.100917
m1038 s44b net09713 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.031397
m1027 net09690 chal44 net09701 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.130524
m1026 vdd! s43a net09690 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.027469
m1025 net09698 net09677 net09701 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.009396
m1024 vdd! s43b net09698 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.139834
m1023 vdd! s43a net09710 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.091202
m1022 net09710 net09681 net09713 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.099353
m1021 vdd! s43b net013342 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.000816
m1020 net013342 chal44 net09713 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.027452
m1019 net09722 chal43 net09733 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.052598
m1018 vdd! s42b net09722 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.051175
m1017 net09730 net09757 net09733 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.008966
m1016 vdd! s42a net09730 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.038943
m1015 vdd! s42b net09742 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.018031
m1014 net09742 net09761 net09745 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.130304
m1013 vdd! s42a net09750 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.101852
m1012 net09750 chal43 net09745 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.120262
m1011 vdd! chal43 net09757 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.128536
m1010 vdd! chal43 net09761 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.058585
m1007 s43b net09733 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.040213
m1006 s43a net09745 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.077666
m995 net09770 chal42 net09781 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.060444
m994 vdd! s41b net09770 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.012866
m993 net09778 net09805 net09781 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.057133
m992 vdd! s41a net09778 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.107885
m991 vdd! s41b net09790 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.079867
m990 net09790 net09809 net09793 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.033696
m989 vdd! s41a net09798 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.002141
m988 net09798 chal42 net09793 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.147912
m985 vdd! chal42 net09805 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.023924
m984 vdd! chal42 net09809 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.001834
m973 s42b net09781 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.050419
m972 s42a net09793 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.016822
m961 vdd! chal41 net09821 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.084449
m960 vdd! chal41 net09825 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.051399
m959 net09826 chal41 net09837 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.000588
m958 vdd! s40a net09826 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.006230
m957 net09834 net09821 net09837 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.053334
m956 vdd! s40b net09834 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.013686
m955 vdd! s40a net09846 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.038357
m954 net09846 net09825 net09849 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.084518
m953 vdd! s40b net09854 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.045583
m952 net09854 chal41 net09849 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.055121
m949 s41a net09837 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.014227
m948 s41b net09849 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.006421
m937 net09866 chal40 net09877 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.006282
m936 vdd! s39b net09866 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.008281
m935 net09874 net09901 net09877 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.014704
m934 vdd! s39a net09874 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.100351
m933 vdd! s39b net09886 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.081243
m932 net09886 net09905 net09889 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.026100
m931 vdd! s39a net09894 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.051781
m930 net09894 chal40 net09889 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.040585
m929 vdd! chal40 net09901 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.050177
m928 vdd! chal40 net09905 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.008558
m925 s40b net09877 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.014509
m924 s40a net09889 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.039583
m921 s39b net09933 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.100745
m920 s39a net09945 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.056024
m909 net09922 chal39 net09933 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.031229
m908 vdd! s38b net09922 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.001607
m907 net09930 net09957 net09933 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.040931
m906 vdd! s38a net09930 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.005837
m905 vdd! s38b net09942 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.001586
m904 net09942 net09961 net09945 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.025024
m903 vdd! s38a net09950 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.038410
m902 net09950 chal39 net09945 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.040354
m901 vdd! chal39 net09957 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.024641
m900 vdd! chal39 net09961 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.042471
m887 net09962 chal38 net09973 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.024693
m886 vdd! s37b net09962 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.106589
m885 net09970 net09985 net09973 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.080319
m884 vdd! s37a net09970 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.072821
m883 s38b net09973 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.136168
m882 vdd! chal38 net09985 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.046299
m881 vdd! chal38 net09989 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.015369
m880 s38a net010001 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.076254
m879 vdd! s37b net09998 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.095070
m878 net09998 net09989 net010001 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.032464
m877 vdd! s37a net010006 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.051497
m876 net010006 chal38 net010001 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.037656
m863 net6849 chal37 net6876 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.050898
m862 vdd! s36a net6849 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.031861
m861 net010018 net010033 net6876 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.068568
m860 vdd! s36b net010018 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.020916
m859 s37a net6876 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.038624
m858 vdd! chal37 net010033 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.013250
m857 vdd! chal37 net5733 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.057105
m856 s37b net010049 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.028919
m855 vdd! s36a net010046 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.034437
m854 net010046 net5733 net010049 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.059632
m853 vdd! s36b net010054 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.154453
m852 net010054 chal37 net010049 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.032939
m851 net010058 chal36 net010069 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.121693
m850 vdd! s35b net010058 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.038876
m849 net010066 net010101 net010069 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.100721
m848 vdd! s35a net010066 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.012929
m847 vdd! s35b net010078 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.056856
m846 net010078 net010105 net010081 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.005785
m845 vdd! s35a net010086 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.028579
m844 net010086 chal36 net010081 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.048609
m833 s36b net010069 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.060150
m832 s36a net010081 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.009058
m1623 vdd! chal69 net12759 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.020144
m819 vdd! chal36 net010101 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.008907
m818 vdd! chal36 net010105 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.020058
m817 s35a net010141 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.029651
m816 s35b net010153 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.103527
m815 s34a net010189 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.023665
m814 s34b net010201 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.066194
m801 vdd! chal35 net010125 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.077954
m800 vdd! chal35 net010129 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.021560
m799 net010130 chal35 net010141 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.060391
m798 vdd! s34a net010130 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.120698
m797 net010138 net010125 net010141 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.023755
m796 vdd! s34b net010138 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.042125
m795 vdd! s34a net010150 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.077820
m794 net010150 net010129 net010153 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.022183
m793 vdd! s34b net010158 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.002610
m792 net010158 chal35 net010153 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.009956
m791 s33b net010229 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.051731
m790 s33a net010241 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.073489
m789 vdd! chal34 net010173 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.032192
m788 vdd! chal34 net010177 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.077708
m783 net010178 chal34 net010189 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.034030
m782 vdd! s33a net010178 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.101915
m781 net010186 net010173 net010189 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.020799
m780 vdd! s33b net010186 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.217189
m779 vdd! s33a net010198 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.012782
m778 net010198 net010177 net010201 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.088198
m777 vdd! s33b net010206 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.022321
m776 net010206 chal34 net010201 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.045545
m775 s32a net010277 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.031419
m774 s32b net010289 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.102480
m773 net010218 chal33 net010229 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.051935
m772 vdd! s32b net010218 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.007930
m771 net010226 net010253 net010229 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.036065
m770 vdd! s32a net010226 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.036283
m769 vdd! s32b net010238 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.012610
m768 net010238 net010257 net010241 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.027832
m767 vdd! s32a net010246 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.000905
m766 net010246 chal33 net010241 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.049103
m765 vdd! chal33 net010253 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.043477
m764 vdd! chal33 net010257 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.099928
m751 vdd! chal32 net010261 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.038285
m750 vdd! chal32 net010265 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.086135
m749 net010266 chal32 net010277 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.006725
m748 vdd! s31a net010266 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.159441
m747 net010274 net010261 net010277 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.008263
m746 vdd! s31b net010274 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.074071
m745 vdd! s31a net010286 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.030541
m744 net010286 net010265 net010289 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.098807
m743 vdd! s31b net010294 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.001023
m742 net010294 chal32 net010289 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.037645
m731 vdd! chal31 net010301 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.128433
m730 vdd! chal31 net010305 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.184487
m729 net010306 chal31 net010317 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.020354
m728 vdd! s30a net010306 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.074592
m727 net010314 net010301 net010317 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.037466
m726 vdd! s30b net010314 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.027114
m725 vdd! s30a net010326 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.022375
m724 net010326 net010305 net010329 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.176717
m723 vdd! s30b net010334 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.070440
m722 net010334 chal31 net010329 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.029691
m711 s31a net010317 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.046284
m710 s31b net010329 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.050930
m707 net010346 chal30 net010357 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.031963
m706 vdd! s29a net010346 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.035432
m705 net010354 net010369 net010357 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.082925
m704 vdd! s29b net010354 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.054725
m703 s30a net010357 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.005627
m702 vdd! chal30 net010369 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.023391
m701 vdd! chal30 net010373 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.024223
m700 s30b net010385 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.008364
m699 vdd! s29a net010382 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.050134
m698 net010382 net010373 net010385 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.015956
m697 vdd! s29b net010390 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.003266
m696 net010390 chal30 net010385 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.074532
m1626 s69a net13861 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.002790
m683 net010394 chal29 net010405 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.064180
m682 vdd! s28b net010394 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.028613
m681 net010402 net5123 net010405 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.028075
m680 vdd! s28a net010402 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.044448
m679 s29b net010405 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.233141
m678 vdd! chal29 net5123 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.050292
m677 vdd! chal29 net010421 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.014278
m676 s29a net6317 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.030094
m675 vdd! s28b net010430 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.107308
m674 net010430 net010421 net6317 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.012859
m673 vdd! s28a net6284 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.022779
m672 net6284 chal29 net6317 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.025372
m659 net010442 chal28 net010453 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.003147
m658 vdd! s27b net010442 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.007167
m657 net010450 net010485 net010453 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.021155
m656 vdd! s27a net010450 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.059752
m655 vdd! s27b net010462 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.050351
m654 net010462 net010489 net010465 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.064192
m653 vdd! s27a net010470 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.048924
m652 net010470 chal28 net010465 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.001811
m641 s28b net010453 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.022964
m640 s28a net010465 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.049074
m627 vdd! chal28 net010485 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.151644
m626 vdd! chal28 net010489 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.003484
m625 s27a net010525 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.043828
m624 s27b net010537 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.080050
m623 s26a net010573 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.127516
m622 s26b net010585 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.020782
m609 vdd! chal27 net010509 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.011096
m608 vdd! chal27 net010513 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.003230
m607 net010514 chal27 net010525 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.007742
m606 vdd! s26a net010514 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.136126
m605 net010522 net010509 net010525 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.081058
m604 vdd! s26b net010522 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.014097
m603 vdd! s26a net010534 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.030925
m602 net010534 net010513 net010537 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.138370
m601 vdd! s26b net010542 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.030716
m600 net010542 chal27 net010537 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.102062
m599 s25b net010613 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.020078
m598 s25a net010625 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.020389
m597 vdd! chal26 net010557 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.101935
m596 vdd! chal26 net010561 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.021214
m591 net010562 chal26 net010573 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.072559
m590 vdd! s25a net010562 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.088019
m589 net010570 net010557 net010573 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.094600
m588 vdd! s25b net010570 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.042029
m587 vdd! s25a net010582 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.006724
m586 net010582 net010561 net010585 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.078452
m585 vdd! s25b net010590 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.039344
m584 net010590 chal26 net010585 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.005758
m583 s24a net010661 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.059050
m582 s24b net010673 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.004263
m581 net010602 chal25 net010613 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.037721
m580 vdd! s24b net010602 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.050525
m579 net010610 net010637 net010613 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.016100
m578 vdd! s24a net010610 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.018909
m577 vdd! s24b net013343 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.092862
m576 net013343 net010641 net010625 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.108929
m575 vdd! s24a net013344 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.130426
m574 net013344 chal25 net010625 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.076612
m573 vdd! chal25 net010637 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.045464
m572 vdd! chal25 net010641 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.091868
m559 vdd! chal24 net013341 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.042447
m558 vdd! chal24 net010649 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.033415
m557 net013345 chal24 net010661 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.021869
m556 vdd! s23a net013345 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.015103
m555 net010658 net013341 net010661 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.094648
m554 vdd! s23b net010658 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.024379
m553 vdd! s23a net010670 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.133511
m552 net010670 net010649 net010673 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.110762
m551 vdd! s23b net010678 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.045058
m550 net010678 chal24 net010673 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.048677
m539 vdd! chal23 net010685 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.046710
m538 vdd! chal23 net013346 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.045809
m537 net010690 chal23 net010701 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.106907
m536 vdd! s22a net010690 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.107210
m535 net010698 net010685 net010701 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.056491
m534 vdd! s22b net010698 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.008377
m533 vdd! s22a net010710 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.074403
m532 net010710 net013346 net010713 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.032754
m531 vdd! s22b net010718 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.204910
m530 net010718 chal23 net010713 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.075959
m519 s23a net010701 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.055700
m518 s23b net010713 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.014547
m515 net010730 chal22 net010741 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.130949
m514 vdd! s21a net010730 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.024257
m513 net010738 net010753 net010741 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.125518
m512 vdd! s21b net010738 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.173787
m511 s22a net010741 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.075107
m510 vdd! chal22 net010753 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.102196
m509 vdd! chal22 net010757 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.015470
m508 s22b net010769 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.003116
m507 vdd! s21a net010766 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.053043
m506 net010766 net010757 net010769 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.126956
m505 vdd! s21b net010774 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.066284
m504 net010774 chal22 net010769 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.019219
m1629 net14388 chal69 net13861 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.038914
m1625 vdd! s68a net14388 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.060000
m491 net010778 chal21 net010789 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.003440
m490 vdd! s20b net010778 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.182404
m489 net010786 net3767 net010789 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.017194
m488 vdd! s20a net010786 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.053853
m487 s21b net010789 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.037897
m486 vdd! chal21 net3767 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.109019
m485 vdd! chal21 net010805 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.078896
m484 s21a net4501 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.037960
m483 vdd! s20b net010814 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.003372
m482 net010814 net010805 net4501 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.003299
m481 vdd! s20a net4447 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.060265
m480 net4447 chal21 net4501 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.145680
m467 s20a net010633 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.067405
m466 s20b net010645 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.023436
m455 s19b net010665 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.021079
m454 s19a net010677 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.065879
m453 vdd! chal20 net010617 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.004928
m452 vdd! chal20 net010621 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.103139
m447 net010622 chal20 net010633 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.086521
m446 vdd! s19a net010622 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.041942
m445 net010630 net010617 net010633 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.108947
m444 vdd! s19b net010630 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.083725
m443 vdd! s19a net010642 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.070626
m442 net010642 net010621 net010645 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.073334
m441 vdd! s19b net010650 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.001815
m440 net010650 chal20 net010645 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.133078
m439 net010654 chal19 net010665 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.008426
m438 vdd! s18b net010654 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.000738
m437 net010662 net010689 net010665 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.015686
m436 vdd! s18a net010662 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.089874
m435 vdd! s18b net010674 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.073767
m434 net010674 net010693 net010677 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.013061
m433 vdd! s18a net010682 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.035018
m432 net010682 chal19 net010677 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.026277
m431 vdd! chal19 net010689 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.025412
m430 vdd! chal19 net010693 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.047686
m409 net4080 chal18 net4091 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.070973
m408 vdd! s17b net4080 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.115152
m407 net4088 net4123 net4091 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.072677
m406 vdd! s17a net4088 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.075456
m405 s18b net4091 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.070423
m404 s18a net4111 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.008852
m403 vdd! s17b net4108 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.049642
m402 net4108 net4127 net4111 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.014059
m401 vdd! s17a net4116 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.010104
m400 net4116 chal18 net4111 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.000137
m387 vdd! chal18 net4123 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.009920
m386 vdd! chal18 net4127 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.009485
m385 s17a net4155 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.031125
m384 s17b net4167 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.086275
m379 vdd! chal17 net4139 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.101295
m378 vdd! chal17 net4143 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.038157
m377 net4144 chal17 net4155 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.004889
m376 vdd! s16a net4144 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.099552
m375 net4152 net4139 net4155 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.025816
m374 vdd! s16b net4152 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.021096
m373 vdd! s16a net4164 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.003974
m372 net4164 net4143 net4167 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.069727
m371 vdd! s16b net4172 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.007131
m370 net4172 chal17 net4167 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.038446
m369 s16b net4195 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.007009
m368 s16a net4207 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.015610
m355 net4184 chal16 net4195 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.138463
m354 vdd! s15b net4184 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.097770
m353 net4192 net4219 net4195 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.070459
m352 vdd! s15a net4192 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.074214
m351 vdd! s15b net4204 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.173240
m350 net4204 net4223 net4207 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.115978
m349 vdd! s15a net4212 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.004135
m348 net4212 chal16 net4207 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.065371
m347 vdd! chal16 net4219 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.041505
m346 vdd! chal16 net4223 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.028956
m345 s15b net4243 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.082155
m344 s15a net4255 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.033320
m333 net4232 chal15 net4243 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.119348
m332 vdd! s14b net4232 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.047577
m331 net4240 net4267 net4243 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.023824
m330 vdd! s14a net4240 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.013575
m329 vdd! s14b net4252 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.015371
m328 net4252 net4271 net4255 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.024025
m327 vdd! s14a net4260 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.039039
m326 net4260 chal15 net4255 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.040001
m325 vdd! chal15 net4267 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.075193
m324 vdd! chal15 net4271 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.076792
m311 net4272 chal14 net4283 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.006575
m310 vdd! s13b net4272 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.031725
m309 net4280 net4295 net4283 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.072438
m308 vdd! s13a net4280 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.080922
m307 s14b net4283 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.079434
m306 vdd! chal14 net4295 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.012339
m305 vdd! chal14 net4299 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.048343
m304 s14a net4311 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.060825
m303 vdd! s13b net4308 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.052608
m302 net4308 net4299 net4311 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.037392
m301 vdd! s13a net4316 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.022001
m300 net4316 chal14 net4311 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.038998
m263 net4320 chal13 net4331 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.048477
m262 vdd! s12a net4320 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.073117
m261 net4328 net4343 net4331 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.121572
m260 vdd! s12b net4328 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.010128
m259 s13a net4331 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.025780
m258 vdd! chal13 net4343 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.119098
m257 vdd! chal13 net4347 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.006525
m256 s13b net4359 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.074721
m255 vdd! s12a net4356 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.106457
m254 net4356 net4347 net4359 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.002958
m253 vdd! s12b net4364 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.040324
m252 net4364 chal13 net4359 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.049487
m1632 net019668 net019691 net13861 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.078561
m1633 vdd! s68b net019668 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.079138
m5 net4368 chal1 net4379 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.090629
m4 vdd! start2 net4368 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.033756
m3 net4376 net4391 net4379 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.095899
m2 vdd! start1 net4376 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.060696
m1 s1b net4379 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.043079
m0 vdd! chal1 net4391 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.008408
m_i_11 vdd! chal1 net4395 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.092523
m_i_1 s1a net4407 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.000477
m_i_7 vdd! start2 net4404 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.014435
m_i_9 net4404 net4395 net4407 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.035465
m_i_8 vdd! start1 net4412 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.063868
m_i_6 net4412 chal1 net4407 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.006392
m24 net4416 chal2 net4427 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.120271
m25 vdd! s1a net4416 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.038600
m26 net4424 net4439 net4427 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.007427
m27 vdd! s1b net4424 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.012432
m28 s2a net4427 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.064227
m29 vdd! chal2 net4439 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.025349
m30 vdd! chal2 net4443 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.014811
m31 s2b net4455 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.166396
m32 vdd! s1a net4452 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.155106
m33 net4452 net4443 net4455 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.096269
m34 vdd! s1b net4460 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.084760
m35 net4460 chal2 net4455 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.060029
m38 vdd! chal3 net4467 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.023959
m39 vdd! chal3 net4471 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.083940
m50 net4472 chal3 net4483 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.032886
m51 vdd! s2a net4472 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.035179
m52 net4480 net4467 net4483 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.133747
m53 vdd! s2b net4480 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.070143
m54 s3a net4483 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.130732
m55 s3b net4503 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.073661
m56 vdd! s2a net4500 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.056255
m57 net4500 net4471 net4503 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.005087
m58 vdd! s2b net4508 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.136640
m59 net4508 chal3 net4503 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.174976
m62 vdd! chal4 net4515 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.084459
m63 vdd! chal4 net4519 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.049519
m74 net4520 chal4 net4531 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.031565
m75 vdd! s3a net4520 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.026279
m76 net4528 net4515 net4531 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.014901
m77 vdd! s3b net4528 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.023049
m78 s4a net4531 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.146445
m79 s4b net4551 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.099524
m80 vdd! s3a net4548 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.067426
m81 net4548 net4519 net4551 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.046018
m82 vdd! s3b net4556 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.075198
m83 net4556 chal4 net4551 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.013921
m84 net4560 chal5 net4571 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.020210
m85 vdd! s4b net4560 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.038212
m86 net4568 net4603 net4571 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.083675
m87 vdd! s4a net4568 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.168356
m88 s5b net4571 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.028948
m89 s5a net4591 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.059035
m90 vdd! s4b net4588 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.059735
m91 net4588 net4607 net4591 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.018378
m92 vdd! s4a net4596 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.100772
m93 net4596 chal5 net4591 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.036735
m104 vdd! chal5 net4603 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.043841
m105 vdd! chal5 net4607 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.034326
m110 vdd! chal6 net4611 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.027449
m111 vdd! chal6 net4615 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.067850
m122 net4616 chal6 net4627 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.004211
m123 vdd! s5a net4616 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.008860
m124 net4624 net4611 net4627 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.040401
m125 vdd! s5b net4624 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.021362
m126 s6a net4627 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.033829
m127 s6b net4647 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.021720
m128 vdd! s5a net4644 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.060308
m129 net4644 net4615 net4647 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.085402
m130 vdd! s5b net4652 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.045185
m131 net4652 chal6 net4647 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.020240
m132 net4656 chal7 net4667 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.070030
m133 vdd! s6b net4656 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.041164
m134 net4664 net4699 net4667 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.109024
m135 vdd! s6a net4664 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.095296
m136 s7b net4667 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.133006
m137 s7a net4687 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.012450
m138 vdd! s6b net4684 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.151663
m139 net4684 net4703 net4687 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.049482
m140 vdd! s6a net4692 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.155773
m141 net4692 chal7 net4687 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.023884
m152 vdd! chal7 net4699 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.157587
m153 vdd! chal7 net4703 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.011630
m156 net4704 chal8 net4715 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.034092
m157 vdd! s7b net4704 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.047108
m158 net4712 net4747 net4715 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.026247
m159 vdd! s7a net4712 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.057434
m160 s8b net4715 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.026241
m161 s8a net4735 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.061494
m162 vdd! s7b net4732 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.069861
m163 net4732 net4751 net4735 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.004932
m164 vdd! s7a net4740 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.020338
m165 net4740 chal8 net4735 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.054484
m176 vdd! chal8 net4747 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.006199
m177 vdd! chal8 net4751 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.103157
m182 vdd! chal9 net4755 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.114786
m183 vdd! chal9 net4759 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.101730
m192 net4760 chal9 net4771 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.056236
m193 vdd! s8a net4760 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.058980
m194 net4768 net4755 net4771 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.003489
m195 vdd! s8b net4768 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.087357
m196 vdd! s8a net4780 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.069097
m197 net4780 net4759 net4783 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.033678
m198 vdd! s8b net4788 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.095256
m199 net4788 chal9 net4783 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.001940
m202 s9a net4771 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.024347
m203 s9b net4783 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.085689
m206 vdd! chal10 net4803 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.051355
m207 vdd! chal10 net4807 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.110569
m208 net4808 chal10 net4819 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.017798
m209 vdd! s9a net4808 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.032507
m210 net4816 net4803 net4819 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.050052
m211 vdd! s9b net4816 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.071109
m212 vdd! s9a net4828 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.012322
m213 net4828 net4807 net4831 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.001491
m214 vdd! s9b net4836 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.102263
m215 net4836 chal10 net4831 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.007731
m226 s10a net4819 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.053806
m227 s10b net4831 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.029495
m230 vdd! chal11 net4851 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.068338
m231 vdd! chal11 net4855 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.132364
m242 net4856 chal11 net4867 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.050794
m243 vdd! s10a net4856 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.018975
m244 net4864 net4851 net4867 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.157610
m245 vdd! s10b net4864 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.181590
m246 s11a net4867 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =-0.118547
m247 s11b net4887 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.062678
m248 vdd! s10a net4884 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.113303
m249 net4884 net4855 net4887 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.044652
m250 vdd! s10b net4892 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.031609
m251 net4892 chal11 net4887 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.012441
m295 s12a net4915 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.057013
m294 s12b net4935 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9 DELVTO =0.061589
m281 net4904 chal12 net4915 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.175417
m280 vdd! s11a net4904 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.033095
m279 net4912 net4923 net4915 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.081759
m278 vdd! s11b net4912 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.162305
m291 vdd! chal12 net4923 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.069850
m290 vdd! chal12 net4927 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =-0.049349
m277 vdd! s11a net4932 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.063501
m276 net4932 net4927 net4935 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.012288
m275 vdd! s11b net4940 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.004777
m274 net4940 chal12 net4935 vdd! PMOS_VTL L=50e-9 W=315e-9 DELVTO =0.000414
xi281 s128a s128b ya yb Arbiter
xi282 clk ya out outb DFF_X1
.param clock_freq=2
.tran 10ps 4ns UIC
.MEASURE TRAN tdlayS1a1 TRIG V(s1a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s1b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS2a1 TRIG V(s2a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s2b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS3a1 TRIG V(s3a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s3b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS4a1 TRIG V(s4a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s4b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS5a1 TRIG V(s5a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s5b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS6a1 TRIG V(s6a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s6b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS7a1 TRIG V(s7a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s7b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS8a1 TRIG V(s8a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s8b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS9a1 TRIG V(s9a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s9b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS10a1 TRIG V(s10a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s10b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS11a1 TRIG V(s11a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s11b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS12a1 TRIG V(s12a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s12b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS13a1 TRIG V(s13a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s13b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS14a1 TRIG V(s14a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s14b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS15a1 TRIG V(s15a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s15b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS16a1 TRIG V(s16a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s16b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS17a1 TRIG V(s17a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s17b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS18a1 TRIG V(s18a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s18b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS19a1 TRIG V(s19a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s19b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS20a1 TRIG V(s20a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s20b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS21a1 TRIG V(s21a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s21b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS22a1 TRIG V(s22a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s22b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS23a1 TRIG V(s23a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s23b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS24a1 TRIG V(s24a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s24b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS25a1 TRIG V(s25a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s25b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS26a1 TRIG V(s26a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s26b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS27a1 TRIG V(s27a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s27b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS28a1 TRIG V(s28a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s28b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS29a1 TRIG V(s29a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s29b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS30a1 TRIG V(s30a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s30b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS31a1 TRIG V(s31a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s31b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS32a1 TRIG V(s32a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s32b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS33a1 TRIG V(s33a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s33b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS34a1 TRIG V(s34a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s34b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS35a1 TRIG V(s35a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s35b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS36a1 TRIG V(s36a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s36b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS37a1 TRIG V(s37a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s37b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS38a1 TRIG V(s38a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s38b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS39a1 TRIG V(s39a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s39b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS40a1 TRIG V(s40a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s40b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS41a1 TRIG V(s41a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s41b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS42a1 TRIG V(s42a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s42b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS43a1 TRIG V(s43a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s43b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS44a1 TRIG V(s44a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s44b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS45a1 TRIG V(s45a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s45b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS46a1 TRIG V(s46a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s46b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS47a1 TRIG V(s47a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s47b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS48a1 TRIG V(s48a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s48b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS49a1 TRIG V(s49a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s49b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS50a1 TRIG V(s50a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s50b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS51a1 TRIG V(s51a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s51b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS52a1 TRIG V(s52a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s52b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS53a1 TRIG V(s53a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s53b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS54a1 TRIG V(s54a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s54b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS55a1 TRIG V(s55a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s55b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS56a1 TRIG V(s56a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s56b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS57a1 TRIG V(s57a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s57b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS58a1 TRIG V(s58a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s58b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS59a1 TRIG V(s59a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s59b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS60a1 TRIG V(s60a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s60b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS61a1 TRIG V(s61a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s61b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS62a1 TRIG V(s62a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s62b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS63a1 TRIG V(s63a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s63b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS64a1 TRIG V(s64a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s64b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS65a1 TRIG V(s65a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s65b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS66a1 TRIG V(s66a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s66b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS67a1 TRIG V(s67a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s67b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS68a1 TRIG V(s68a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s68b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS69a1 TRIG V(s69a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s69b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS70a1 TRIG V(s70a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s70b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS71a1 TRIG V(s71a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s71b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS72a1 TRIG V(s72a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s72b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS73a1 TRIG V(s73a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s73b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS74a1 TRIG V(s74a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s74b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS75a1 TRIG V(s75a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s75b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS76a1 TRIG V(s76a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s76b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS77a1 TRIG V(s77a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s77b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS78a1 TRIG V(s78a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s78b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS79a1 TRIG V(s79a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s79b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS80a1 TRIG V(s80a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s80b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS81a1 TRIG V(s81a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s81b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS82a1 TRIG V(s82a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s82b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS83a1 TRIG V(s83a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s83b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS84a1 TRIG V(s84a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s84b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS85a1 TRIG V(s85a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s85b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS86a1 TRIG V(s86a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s86b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS87a1 TRIG V(s87a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s87b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS88a1 TRIG V(s88a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s88b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS89a1 TRIG V(s89a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s89b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS90a1 TRIG V(s90a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s90b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS91a1 TRIG V(s91a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s91b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS92a1 TRIG V(s92a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s92b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS93a1 TRIG V(s93a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s93b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS94a1 TRIG V(s94a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s94b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS95a1 TRIG V(s95a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s95b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS96a1 TRIG V(s96a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s96b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS97a1 TRIG V(s97a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s97b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS98a1 TRIG V(s98a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s98b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS99a1 TRIG V(s99a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s99b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS100a1 TRIG V(s100a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s100b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS101a1 TRIG V(s101a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s101b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS102a1 TRIG V(s102a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s102b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS103a1 TRIG V(s103a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s103b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS104a1 TRIG V(s104a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s104b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS105a1 TRIG V(s105a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s105b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS106a1 TRIG V(s106a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s106b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS107a1 TRIG V(s107a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s107b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS108a1 TRIG V(s108a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s108b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS109a1 TRIG V(s109a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s109b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS110a1 TRIG V(s110a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s110b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS111a1 TRIG V(s111a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s111b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS112a1 TRIG V(s112a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s112b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS113a1 TRIG V(s113a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s113b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS114a1 TRIG V(s114a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s114b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS115a1 TRIG V(s115a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s115b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS116a1 TRIG V(s116a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s116b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS117a1 TRIG V(s117a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s117b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS118a1 TRIG V(s118a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s118b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS119a1 TRIG V(s119a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s119b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS120a1 TRIG V(s120a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s120b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS121a1 TRIG V(s121a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s121b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS122a1 TRIG V(s122a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s122b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS123a1 TRIG V(s123a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s123b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS124a1 TRIG V(s124a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s124b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS125a1 TRIG V(s125a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s125b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS126a1 TRIG V(s126a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s126b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS127a1 TRIG V(s127a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s127b) VAL = 0.5 RISE = 1
.MEASURE TRAN tdlayS128a1 TRIG V(s128a) VAL = 0.5 RISE = 1 TD=0.5ns TARG V(s128b) VAL = 0.5 RISE = 1
.MEASURE TRAN PowEva1 INTEG I(vsupply) From=0.52ns TO=3.99ns
.MEASURE TRAN PowEva3Half1 INTEG I(vsupply) From=3.25ns TO=3.75ns
.MEASURE TRAN ya1 AVG V(ya) FROM=3.991ns TO=3.9911ns
.MEASURE TRAN outa1 AVG V(out) FROM=3.991ns TO=3.9911ns
.IC I(vsupply)=0 V(start1)=0 V(start2)=0 V(ya)=0 V(out)=0
.PRINT TRAN I(vsupply)
.END
